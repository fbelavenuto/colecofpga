-- generated with romgen v3.0 by MikeJ
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity biosx is
	port (
		CLK		: in    std_logic;
		ENA		: in    std_logic;
		ADDR		: in    std_logic_vector(12 downto 0);
		DATA		: out   std_logic_vector(7 downto 0)
	);
end;

architecture RTL of biosx is

  type ROM_ARRAY is array(0 to 8191) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"31",x"B9",x"73",x"C3",x"6E",x"00",x"FF",x"FF", -- 0x0000
    x"C3",x"0C",x"80",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0008
    x"C3",x"0F",x"80",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0010
    x"C3",x"12",x"80",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0018
    x"C3",x"15",x"80",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0020
    x"C3",x"18",x"80",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0028
    x"C3",x"1B",x"80",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0030
    x"C3",x"1E",x"80",x"2A",x"C8",x"73",x"CB",x"7C", -- 0x0038
    x"28",x"06",x"CB",x"44",x"28",x"06",x"18",x"07", -- 0x0040
    x"CB",x"44",x"28",x"03",x"37",x"18",x"01",x"B7", -- 0x0048
    x"CB",x"15",x"CB",x"14",x"22",x"C8",x"73",x"7D", -- 0x0050
    x"C9",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0058
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"C3",x"21", -- 0x0060
    x"80",x"3C",x"AB",x"16",x"23",x"16",x"2A",x"00", -- 0x0068
    x"80",x"7D",x"FE",x"55",x"C2",x"81",x"00",x"7C", -- 0x0070
    x"FE",x"AA",x"C2",x"81",x"00",x"2A",x"0A",x"80", -- 0x0078
    x"E9",x"CD",x"D6",x"1F",x"21",x"33",x"00",x"22", -- 0x0080
    x"C8",x"73",x"CD",x"05",x"11",x"3E",x"00",x"32", -- 0x0088
    x"C6",x"73",x"32",x"C7",x"73",x"C3",x"19",x"13", -- 0x0090
    x"E1",x"E3",x"E5",x"0A",x"6F",x"03",x"0A",x"03", -- 0x0098
    x"67",x"E3",x"D5",x"5E",x"23",x"56",x"23",x"E5", -- 0x00A0
    x"7B",x"B2",x"C2",x"B7",x"00",x"E1",x"5E",x"23", -- 0x00A8
    x"56",x"23",x"E5",x"EB",x"5E",x"23",x"56",x"03", -- 0x00B0
    x"0A",x"07",x"D2",x"DA",x"00",x"03",x"E1",x"E3", -- 0x00B8
    x"73",x"23",x"72",x"23",x"D1",x"E3",x"2B",x"AF", -- 0x00C0
    x"BC",x"C2",x"D0",x"00",x"BD",x"CA",x"D6",x"00", -- 0x00C8
    x"E3",x"E5",x"EB",x"C3",x"A3",x"00",x"E1",x"EB", -- 0x00D0
    x"E3",x"E9",x"E1",x"E3",x"E5",x"0F",x"67",x"0B", -- 0x00D8
    x"0A",x"6F",x"E3",x"03",x"03",x"1A",x"77",x"23", -- 0x00E0
    x"13",x"E3",x"2B",x"AF",x"BD",x"C2",x"F4",x"00", -- 0x00E8
    x"BC",x"CA",x"F8",x"00",x"E3",x"C3",x"E5",x"00", -- 0x00F0
    x"E1",x"C3",x"C4",x"00",x"DD",x"7E",x"07",x"FE", -- 0x00F8
    x"00",x"20",x"09",x"DD",x"7E",x"05",x"3D",x"C8", -- 0x0100
    x"DD",x"77",x"05",x"C9",x"DD",x"E5",x"E1",x"1E", -- 0x0108
    x"06",x"16",x"00",x"19",x"CD",x"90",x"01",x"20", -- 0x0110
    x"15",x"CD",x"A6",x"01",x"2B",x"7E",x"3D",x"C8", -- 0x0118
    x"77",x"2B",x"2B",x"DD",x"7E",x"07",x"CD",x"B1", -- 0x0120
    x"01",x"23",x"CB",x"96",x"F6",x"FF",x"C9",x"DD", -- 0x0128
    x"7E",x"08",x"FE",x"00",x"C8",x"DD",x"E5",x"E1", -- 0x0130
    x"16",x"00",x"1E",x"09",x"19",x"CD",x"90",x"01", -- 0x0138
    x"20",x"21",x"CD",x"A6",x"01",x"2B",x"CD",x"90", -- 0x0140
    x"01",x"28",x"16",x"7E",x"E6",x"F0",x"5F",x"2B", -- 0x0148
    x"2B",x"2B",x"2B",x"7E",x"E6",x"F0",x"83",x"5F", -- 0x0150
    x"7E",x"E6",x"0F",x"B3",x"77",x"F6",x"FF",x"18", -- 0x0158
    x"02",x"36",x"00",x"C9",x"DD",x"7E",x"04",x"CB", -- 0x0160
    x"61",x"28",x"04",x"0F",x"0F",x"0F",x"0F",x"E6", -- 0x0168
    x"0F",x"B1",x"D3",x"FF",x"C9",x"DD",x"7E",x"03", -- 0x0170
    x"E6",x"0F",x"B2",x"D3",x"FF",x"DD",x"7E",x"03", -- 0x0178
    x"E6",x"F0",x"57",x"DD",x"7E",x"04",x"E6",x"0F", -- 0x0180
    x"B2",x"0F",x"0F",x"0F",x"0F",x"D3",x"FF",x"C9", -- 0x0188
    x"3E",x"00",x"ED",x"67",x"D6",x"01",x"F5",x"ED", -- 0x0190
    x"6F",x"F1",x"C9",x"3E",x"00",x"ED",x"6F",x"D6", -- 0x0198
    x"01",x"F5",x"ED",x"67",x"F1",x"C9",x"7E",x"E6", -- 0x01A0
    x"F0",x"47",x"0F",x"0F",x"0F",x"0F",x"B0",x"77", -- 0x01A8
    x"C9",x"06",x"00",x"CB",x"7F",x"28",x"02",x"06", -- 0x01B0
    x"FF",x"86",x"77",x"23",x"7E",x"88",x"77",x"2B", -- 0x01B8
    x"C9",x"2A",x"20",x"70",x"2B",x"2B",x"48",x"06", -- 0x01C0
    x"00",x"CB",x"01",x"CB",x"01",x"09",x"5E",x"23", -- 0x01C8
    x"56",x"D5",x"DD",x"E1",x"C9",x"DD",x"75",x"01", -- 0x01D0
    x"DD",x"74",x"02",x"1A",x"E6",x"3F",x"47",x"DD", -- 0x01D8
    x"7E",x"00",x"E6",x"C0",x"B0",x"DD",x"77",x"00", -- 0x01E0
    x"C9",x"DD",x"7E",x"00",x"FE",x"FF",x"C8",x"E6", -- 0x01E8
    x"3F",x"FE",x"3E",x"C0",x"DD",x"E5",x"E1",x"23", -- 0x01F0
    x"5E",x"23",x"56",x"EB",x"C9",x"02",x"00",x"01", -- 0x01F8
    x"00",x"02",x"00",x"01",x"FD",x"01",x"11",x"BA", -- 0x0200
    x"73",x"CD",x"98",x"00",x"3A",x"BA",x"73",x"47", -- 0x0208
    x"2A",x"BB",x"73",x"22",x"20",x"70",x"23",x"23", -- 0x0210
    x"5E",x"23",x"56",x"EB",x"1E",x"0A",x"16",x"00", -- 0x0218
    x"36",x"FF",x"19",x"10",x"FB",x"36",x"00",x"21", -- 0x0220
    x"4C",x"02",x"22",x"22",x"70",x"22",x"24",x"70", -- 0x0228
    x"22",x"26",x"70",x"22",x"28",x"70",x"3E",x"FF", -- 0x0230
    x"32",x"2A",x"70",x"3E",x"9F",x"D3",x"FF",x"3E", -- 0x0238
    x"BF",x"D3",x"FF",x"3E",x"DF",x"D3",x"FF",x"3E", -- 0x0240
    x"FF",x"D3",x"FF",x"C9",x"FF",x"01",x"00",x"01", -- 0x0248
    x"00",x"01",x"4D",x"02",x"11",x"BA",x"73",x"CD", -- 0x0250
    x"98",x"00",x"3A",x"BA",x"73",x"47",x"C5",x"CD", -- 0x0258
    x"C1",x"01",x"DD",x"7E",x"00",x"E6",x"3F",x"C1", -- 0x0260
    x"B8",x"C8",x"DD",x"70",x"00",x"2B",x"2B",x"56", -- 0x0268
    x"2B",x"5E",x"DD",x"73",x"01",x"DD",x"72",x"02", -- 0x0270
    x"CD",x"5F",x"03",x"CD",x"95",x"02",x"C9",x"06", -- 0x0278
    x"01",x"CD",x"C1",x"01",x"3E",x"00",x"DD",x"BE", -- 0x0280
    x"00",x"C8",x"CD",x"D6",x"02",x"1E",x"0A",x"16", -- 0x0288
    x"00",x"DD",x"19",x"18",x"EF",x"DD",x"E5",x"21", -- 0x0290
    x"4C",x"02",x"22",x"22",x"70",x"22",x"24",x"70", -- 0x0298
    x"22",x"26",x"70",x"22",x"28",x"70",x"06",x"01", -- 0x02A0
    x"CD",x"C1",x"01",x"DD",x"7E",x"00",x"FE",x"00", -- 0x02A8
    x"28",x"21",x"FE",x"FF",x"28",x"15",x"DD",x"7E", -- 0x02B0
    x"00",x"E6",x"C0",x"07",x"07",x"07",x"5F",x"16", -- 0x02B8
    x"00",x"21",x"22",x"70",x"19",x"DD",x"E5",x"D1", -- 0x02C0
    x"73",x"23",x"72",x"1E",x"0A",x"16",x"00",x"DD", -- 0x02C8
    x"19",x"18",x"D8",x"DD",x"E1",x"C9",x"CD",x"E9", -- 0x02D0
    x"01",x"FE",x"FF",x"C8",x"FE",x"3E",x"20",x"06", -- 0x02D8
    x"1E",x"07",x"16",x"00",x"19",x"E9",x"CD",x"2F", -- 0x02E0
    x"01",x"CD",x"FC",x"00",x"20",x"11",x"DD",x"7E", -- 0x02E8
    x"00",x"F5",x"CD",x"5F",x"03",x"C1",x"DD",x"7E", -- 0x02F0
    x"00",x"B8",x"28",x"03",x"CD",x"95",x"02",x"C9", -- 0x02F8
    x"3E",x"9F",x"0E",x"90",x"16",x"80",x"DD",x"2A", -- 0x0300
    x"24",x"70",x"CD",x"4E",x"03",x"3E",x"BF",x"0E", -- 0x0308
    x"B0",x"16",x"A0",x"DD",x"2A",x"26",x"70",x"CD", -- 0x0310
    x"4E",x"03",x"3E",x"DF",x"0E",x"D0",x"16",x"C0", -- 0x0318
    x"DD",x"2A",x"28",x"70",x"CD",x"4E",x"03",x"3E", -- 0x0320
    x"FF",x"0E",x"F0",x"DD",x"2A",x"22",x"70",x"DD", -- 0x0328
    x"5E",x"00",x"1C",x"20",x"04",x"D3",x"FF",x"18", -- 0x0330
    x"14",x"CD",x"64",x"01",x"DD",x"7E",x"04",x"E6", -- 0x0338
    x"0F",x"21",x"2A",x"70",x"BE",x"28",x"06",x"77", -- 0x0340
    x"0E",x"E0",x"CD",x"64",x"01",x"C9",x"DD",x"5E", -- 0x0348
    x"00",x"1C",x"20",x"04",x"D3",x"FF",x"18",x"06", -- 0x0350
    x"CD",x"64",x"01",x"CD",x"75",x"01",x"C9",x"DD", -- 0x0358
    x"7E",x"00",x"E6",x"3F",x"F5",x"DD",x"36",x"00", -- 0x0360
    x"FF",x"DD",x"6E",x"01",x"DD",x"66",x"02",x"7E", -- 0x0368
    x"47",x"CB",x"6F",x"28",x"1C",x"C5",x"E6",x"1F", -- 0x0370
    x"23",x"DD",x"75",x"01",x"DD",x"74",x"02",x"DD", -- 0x0378
    x"36",x"04",x"F0",x"DD",x"77",x"05",x"DD",x"36", -- 0x0380
    x"07",x"00",x"DD",x"36",x"08",x"00",x"C3",x"61", -- 0x0388
    x"04",x"CB",x"67",x"28",x"0F",x"CB",x"5F",x"28", -- 0x0390
    x"05",x"C1",x"CD",x"5E",x"02",x"C9",x"3E",x"FF", -- 0x0398
    x"F5",x"C3",x"61",x"04",x"E6",x"3C",x"FE",x"04", -- 0x03A0
    x"20",x"28",x"FD",x"E1",x"FD",x"E5",x"C5",x"23", -- 0x03A8
    x"5E",x"DD",x"73",x"01",x"23",x"56",x"DD",x"72", -- 0x03B0
    x"02",x"23",x"FD",x"E5",x"F1",x"D5",x"FD",x"E1", -- 0x03B8
    x"11",x"C6",x"03",x"D5",x"FD",x"E9",x"16",x"00", -- 0x03C0
    x"1E",x"07",x"FD",x"19",x"11",x"61",x"04",x"D5", -- 0x03C8
    x"FD",x"E9",x"C5",x"78",x"E6",x"03",x"FE",x"00", -- 0x03D0
    x"20",x"20",x"23",x"23",x"23",x"23",x"DD",x"75", -- 0x03D8
    x"01",x"DD",x"74",x"02",x"2B",x"11",x"05",x"00", -- 0x03E0
    x"CD",x"78",x"04",x"01",x"03",x"00",x"ED",x"B8", -- 0x03E8
    x"DD",x"36",x"07",x"00",x"DD",x"36",x"08",x"00", -- 0x03F0
    x"18",x"67",x"FE",x"01",x"20",x"1B",x"1E",x"06", -- 0x03F8
    x"16",x"00",x"19",x"DD",x"75",x"01",x"DD",x"74", -- 0x0400
    x"02",x"2B",x"1C",x"CD",x"78",x"04",x"01",x"05", -- 0x0408
    x"00",x"ED",x"B8",x"DD",x"36",x"08",x"00",x"18", -- 0x0410
    x"48",x"FE",x"02",x"20",x"28",x"1E",x"06",x"16", -- 0x0418
    x"00",x"19",x"F1",x"F5",x"E6",x"C0",x"20",x"01", -- 0x0420
    x"2B",x"DD",x"75",x"01",x"DD",x"74",x"02",x"2B", -- 0x0428
    x"1E",x"09",x"CD",x"78",x"04",x"01",x"02",x"00", -- 0x0430
    x"ED",x"B8",x"3E",x"00",x"12",x"1B",x"1B",x"0E", -- 0x0438
    x"03",x"ED",x"B8",x"18",x"1C",x"1E",x"08",x"16", -- 0x0440
    x"00",x"19",x"DD",x"75",x"01",x"DD",x"74",x"02", -- 0x0448
    x"2B",x"DD",x"E5",x"FD",x"E1",x"1E",x"09",x"FD", -- 0x0450
    x"19",x"FD",x"E5",x"D1",x"01",x"07",x"00",x"ED", -- 0x0458
    x"B8",x"DD",x"E5",x"E1",x"F1",x"C1",x"FE",x"FF", -- 0x0460
    x"C8",x"57",x"E6",x"3F",x"FE",x"04",x"20",x"02", -- 0x0468
    x"06",x"3E",x"7A",x"E6",x"C0",x"B0",x"77",x"C9", -- 0x0470
    x"DD",x"E5",x"FD",x"E1",x"FD",x"19",x"FD",x"E5", -- 0x0478
    x"D1",x"C9",x"02",x"00",x"FE",x"FF",x"01",x"00", -- 0x0480
    x"01",x"82",x"04",x"11",x"BA",x"73",x"CD",x"98", -- 0x0488
    x"00",x"2A",x"BA",x"73",x"5E",x"23",x"56",x"EB", -- 0x0490
    x"3A",x"BC",x"73",x"FE",x"00",x"28",x"03",x"37", -- 0x0498
    x"18",x"01",x"B7",x"5E",x"23",x"56",x"23",x"4E", -- 0x04A0
    x"23",x"46",x"23",x"3E",x"00",x"02",x"1A",x"F5", -- 0x04A8
    x"E6",x"0F",x"CA",x"E7",x"04",x"3D",x"CA",x"F1", -- 0x04B0
    x"05",x"3D",x"CA",x"00",x"06",x"3D",x"CA",x"00", -- 0x04B8
    x"06",x"3D",x"28",x"02",x"F1",x"C9",x"1A",x"1F", -- 0x04C0
    x"1F",x"1F",x"1F",x"E6",x"0F",x"47",x"5E",x"23", -- 0x04C8
    x"56",x"23",x"B7",x"28",x"10",x"F1",x"F5",x"E5", -- 0x04D0
    x"C5",x"EB",x"CD",x"A3",x"04",x"C1",x"E1",x"5E", -- 0x04D8
    x"23",x"56",x"23",x"10",x"F0",x"F1",x"C9",x"CD", -- 0x04E0
    x"72",x"05",x"1A",x"6F",x"13",x"1A",x"85",x"FD", -- 0x04E8
    x"77",x"05",x"26",x"00",x"F1",x"30",x"38",x"F5", -- 0x04F0
    x"3A",x"C3",x"73",x"CB",x"4F",x"28",x"31",x"EB", -- 0x04F8
    x"44",x"4D",x"6E",x"26",x"00",x"E5",x"29",x"29", -- 0x0500
    x"29",x"E5",x"03",x"0A",x"6F",x"03",x"0A",x"67", -- 0x0508
    x"C1",x"FD",x"E1",x"F1",x"CB",x"7F",x"28",x"03", -- 0x0510
    x"CD",x"94",x"05",x"CD",x"E8",x"05",x"CB",x"77", -- 0x0518
    x"28",x"03",x"CD",x"94",x"05",x"CD",x"E8",x"05", -- 0x0520
    x"CB",x"6F",x"28",x"03",x"CD",x"94",x"05",x"C9", -- 0x0528
    x"EB",x"4E",x"06",x"00",x"C5",x"FD",x"E1",x"23", -- 0x0530
    x"7E",x"23",x"66",x"6F",x"E5",x"C5",x"D5",x"FD", -- 0x0538
    x"E5",x"3E",x"03",x"CD",x"27",x"1C",x"C1",x"E1", -- 0x0540
    x"5D",x"54",x"09",x"2B",x"CB",x"3C",x"CB",x"1D", -- 0x0548
    x"CB",x"3C",x"CB",x"1D",x"CB",x"3C",x"CB",x"1D", -- 0x0550
    x"CB",x"2B",x"CB",x"2B",x"CB",x"2B",x"B7",x"ED", -- 0x0558
    x"52",x"23",x"E5",x"FD",x"E1",x"E1",x"29",x"29", -- 0x0560
    x"29",x"C1",x"09",x"3E",x"04",x"CD",x"27",x"1C", -- 0x0568
    x"F1",x"C9",x"C5",x"FD",x"E1",x"D5",x"5E",x"23", -- 0x0570
    x"56",x"CB",x"7A",x"20",x"14",x"7A",x"FE",x"70", -- 0x0578
    x"38",x"06",x"3E",x"80",x"12",x"18",x"0A",x"80", -- 0x0580
    x"21",x"87",x"05",x"01",x"01",x"00",x"CD",x"01", -- 0x0588
    x"1D",x"D1",x"13",x"C9",x"F5",x"C5",x"FD",x"E5", -- 0x0590
    x"D5",x"E5",x"3E",x"03",x"CD",x"27",x"1C",x"E1", -- 0x0598
    x"D1",x"FD",x"E1",x"C1",x"F1",x"F5",x"C5",x"FD", -- 0x05A0
    x"E5",x"D5",x"E5",x"CB",x"67",x"20",x"0D",x"09", -- 0x05A8
    x"3E",x"04",x"CD",x"27",x"1C",x"E1",x"D1",x"FD", -- 0x05B0
    x"E1",x"C1",x"F1",x"C9",x"09",x"4D",x"44",x"FD", -- 0x05B8
    x"E5",x"E1",x"E5",x"0A",x"C5",x"01",x"08",x"00", -- 0x05C0
    x"2A",x"06",x"80",x"09",x"06",x"08",x"2B",x"77", -- 0x05C8
    x"10",x"FC",x"D5",x"FD",x"21",x"01",x"00",x"3E", -- 0x05D0
    x"04",x"CD",x"27",x"1C",x"D1",x"C1",x"13",x"03", -- 0x05D8
    x"E1",x"2B",x"7C",x"B5",x"20",x"DC",x"18",x"CD", -- 0x05E0
    x"C5",x"01",x"00",x"01",x"EB",x"09",x"EB",x"C1", -- 0x05E8
    x"C9",x"CD",x"72",x"05",x"13",x"1A",x"FD",x"77", -- 0x05F0
    x"05",x"13",x"1A",x"FD",x"77",x"06",x"F1",x"C9", -- 0x05F8
    x"03",x"03",x"03",x"03",x"03",x"EB",x"23",x"7E", -- 0x0600
    x"5F",x"16",x"00",x"D5",x"23",x"5E",x"23",x"56", -- 0x0608
    x"23",x"86",x"02",x"4E",x"06",x"00",x"C5",x"FD", -- 0x0610
    x"E1",x"EB",x"D1",x"F1",x"D0",x"3E",x"01",x"CD", -- 0x0618
    x"27",x"1C",x"C9",x"DD",x"E5",x"2A",x"CD",x"73", -- 0x0620
    x"D1",x"73",x"23",x"72",x"23",x"70",x"23",x"EB", -- 0x0628
    x"3A",x"CB",x"73",x"3C",x"21",x"CA",x"73",x"BE", -- 0x0630
    x"20",x"0D",x"3E",x"00",x"32",x"CB",x"73",x"2A", -- 0x0638
    x"D1",x"73",x"22",x"CD",x"73",x"18",x"07",x"32", -- 0x0640
    x"CB",x"73",x"ED",x"53",x"CD",x"73",x"C9",x"02", -- 0x0648
    x"00",x"01",x"00",x"FE",x"FF",x"01",x"4F",x"06", -- 0x0650
    x"11",x"BA",x"73",x"CD",x"98",x"00",x"3A",x"BA", -- 0x0658
    x"73",x"2A",x"BB",x"73",x"32",x"CA",x"73",x"3E", -- 0x0660
    x"00",x"32",x"CB",x"73",x"32",x"CC",x"73",x"22", -- 0x0668
    x"D1",x"73",x"22",x"CD",x"73",x"22",x"CF",x"73", -- 0x0670
    x"C9",x"3A",x"C6",x"73",x"F5",x"3E",x"00",x"32", -- 0x0678
    x"C6",x"73",x"3A",x"CC",x"73",x"21",x"CB",x"73", -- 0x0680
    x"BE",x"28",x"31",x"2A",x"CF",x"73",x"5E",x"23", -- 0x0688
    x"56",x"23",x"46",x"23",x"D5",x"DD",x"E1",x"E5", -- 0x0690
    x"CD",x"E3",x"06",x"3A",x"CC",x"73",x"3C",x"21", -- 0x0698
    x"CA",x"73",x"BE",x"20",x"0E",x"3E",x"00",x"32", -- 0x06A0
    x"CC",x"73",x"2A",x"D1",x"73",x"22",x"CF",x"73", -- 0x06A8
    x"E1",x"18",x"07",x"32",x"CC",x"73",x"E1",x"22", -- 0x06B0
    x"CF",x"73",x"18",x"C6",x"F1",x"32",x"C6",x"73", -- 0x06B8
    x"C9",x"02",x"00",x"02",x"00",x"01",x"00",x"01", -- 0x06C0
    x"C1",x"06",x"11",x"BA",x"73",x"CD",x"98",x"00", -- 0x06C8
    x"DD",x"2A",x"BA",x"73",x"3A",x"BC",x"73",x"47", -- 0x06D0
    x"3A",x"C6",x"73",x"FE",x"01",x"20",x"04",x"CD", -- 0x06D8
    x"23",x"06",x"C9",x"DD",x"66",x"01",x"DD",x"6E", -- 0x06E0
    x"00",x"7E",x"4F",x"E6",x"0F",x"CA",x"FF",x"06", -- 0x06E8
    x"3D",x"CA",x"87",x"0A",x"3D",x"CA",x"DF",x"08", -- 0x06F0
    x"3D",x"CA",x"55",x"09",x"C3",x"A2",x"0E",x"DD", -- 0x06F8
    x"56",x"03",x"DD",x"5E",x"02",x"D5",x"FD",x"E1", -- 0x0700
    x"FD",x"56",x"02",x"FD",x"5E",x"01",x"CD",x"E8", -- 0x0708
    x"07",x"4B",x"FD",x"56",x"04",x"FD",x"5E",x"03", -- 0x0710
    x"CD",x"E8",x"07",x"43",x"FD",x"5E",x"00",x"16", -- 0x0718
    x"00",x"19",x"19",x"1E",x"05",x"19",x"5E",x"23", -- 0x0720
    x"56",x"EB",x"C5",x"D1",x"4E",x"23",x"46",x"23", -- 0x0728
    x"DD",x"7E",x"05",x"CB",x"7F",x"28",x"04",x"CD", -- 0x0730
    x"0B",x"08",x"C9",x"C5",x"D5",x"E5",x"FE",x"70", -- 0x0738
    x"28",x"02",x"38",x"07",x"67",x"DD",x"6E",x"04", -- 0x0740
    x"7E",x"18",x"35",x"2A",x"06",x"80",x"DD",x"56", -- 0x0748
    x"05",x"DD",x"5E",x"04",x"E5",x"D5",x"E5",x"01", -- 0x0750
    x"04",x"00",x"CD",x"3E",x"1D",x"E1",x"7E",x"FE", -- 0x0758
    x"80",x"20",x"03",x"D1",x"18",x"19",x"23",x"23", -- 0x0760
    x"46",x"23",x"5E",x"16",x"00",x"23",x"EB",x"18", -- 0x0768
    x"01",x"29",x"10",x"FD",x"E5",x"C1",x"EB",x"D1", -- 0x0770
    x"13",x"13",x"13",x"13",x"CD",x"3E",x"1D",x"E1", -- 0x0778
    x"7E",x"FE",x"80",x"28",x"0F",x"5E",x"23",x"56", -- 0x0780
    x"23",x"4E",x"23",x"46",x"23",x"DD",x"E5",x"CD", -- 0x0788
    x"0B",x"08",x"DD",x"E1",x"E1",x"D1",x"C1",x"C5", -- 0x0790
    x"D5",x"E5",x"DD",x"66",x"05",x"DD",x"6E",x"04", -- 0x0798
    x"3E",x"70",x"BC",x"38",x"03",x"2A",x"06",x"80", -- 0x07A0
    x"73",x"23",x"72",x"23",x"71",x"23",x"70",x"23", -- 0x07A8
    x"DD",x"E5",x"CD",x"98",x"08",x"DD",x"E1",x"E1", -- 0x07B0
    x"D1",x"C1",x"DD",x"E5",x"CD",x"0B",x"08",x"DD", -- 0x07B8
    x"E1",x"DD",x"56",x"05",x"3E",x"70",x"BA",x"28", -- 0x07C0
    x"1E",x"38",x"1C",x"DD",x"5E",x"04",x"D9",x"2A", -- 0x07C8
    x"06",x"80",x"E5",x"23",x"23",x"5E",x"16",x"00", -- 0x07D0
    x"23",x"46",x"EB",x"18",x"01",x"29",x"10",x"FD", -- 0x07D8
    x"E5",x"D9",x"C1",x"E1",x"CD",x"01",x"1D",x"C9", -- 0x07E0
    x"E5",x"CB",x"2A",x"CB",x"1B",x"CB",x"2A",x"CB", -- 0x07E8
    x"1B",x"CB",x"2A",x"CB",x"1B",x"CB",x"7A",x"20", -- 0x07F0
    x"09",x"21",x"80",x"FF",x"19",x"E1",x"D0",x"1E", -- 0x07F8
    x"7F",x"C9",x"21",x"80",x"00",x"19",x"E1",x"D8", -- 0x0800
    x"1E",x"80",x"C9",x"C5",x"D5",x"E5",x"D9",x"E1", -- 0x0808
    x"D1",x"C1",x"CD",x"C0",x"08",x"D9",x"7B",x"CB", -- 0x0810
    x"7F",x"20",x"03",x"FE",x"20",x"D0",x"81",x"CB", -- 0x0818
    x"7F",x"C0",x"B7",x"C8",x"CB",x"7B",x"28",x"20", -- 0x0820
    x"79",x"83",x"D5",x"FE",x"21",x"38",x"02",x"3E", -- 0x0828
    x"20",x"5F",x"16",x"00",x"D5",x"FD",x"E1",x"D1", -- 0x0830
    x"7B",x"D9",x"C5",x"ED",x"44",x"4F",x"06",x"00", -- 0x0838
    x"09",x"EB",x"09",x"EB",x"C1",x"D9",x"18",x"1C", -- 0x0840
    x"7B",x"81",x"FE",x"1F",x"28",x"0F",x"38",x"0D", -- 0x0848
    x"3E",x"20",x"93",x"D5",x"5F",x"16",x"00",x"D5", -- 0x0850
    x"FD",x"E1",x"D1",x"18",x"07",x"C5",x"06",x"00", -- 0x0858
    x"C5",x"FD",x"E1",x"C1",x"1E",x"00",x"7A",x"83", -- 0x0860
    x"CB",x"7F",x"20",x"19",x"FE",x"18",x"30",x"15", -- 0x0868
    x"C5",x"D5",x"D9",x"C5",x"D5",x"E5",x"FD",x"E5", -- 0x0870
    x"3E",x"02",x"CD",x"27",x"1C",x"FD",x"E1",x"E1", -- 0x0878
    x"D1",x"C1",x"D9",x"D1",x"C1",x"D9",x"C5",x"06", -- 0x0880
    x"00",x"09",x"EB",x"01",x"20",x"00",x"09",x"EB", -- 0x0888
    x"C1",x"D9",x"1C",x"7B",x"B8",x"20",x"CF",x"C9", -- 0x0890
    x"CD",x"C0",x"08",x"C5",x"06",x"00",x"C5",x"FD", -- 0x0898
    x"E1",x"C1",x"C5",x"D5",x"E5",x"FD",x"E5",x"3E", -- 0x08A0
    x"02",x"CD",x"A3",x"1B",x"FD",x"E1",x"E1",x"D1", -- 0x08A8
    x"C1",x"C5",x"06",x"00",x"09",x"01",x"20",x"00", -- 0x08B0
    x"EB",x"09",x"EB",x"C1",x"05",x"20",x"E3",x"C9", -- 0x08B8
    x"E5",x"CB",x"7A",x"28",x"04",x"26",x"FF",x"18", -- 0x08C0
    x"02",x"26",x"00",x"6A",x"29",x"29",x"29",x"29", -- 0x08C8
    x"29",x"CB",x"7B",x"28",x"04",x"16",x"FF",x"18", -- 0x08D0
    x"02",x"16",x"00",x"19",x"EB",x"E1",x"C9",x"FD", -- 0x08D8
    x"2A",x"06",x"80",x"DD",x"6E",x"02",x"DD",x"66", -- 0x08E0
    x"03",x"11",x"01",x"00",x"19",x"4E",x"23",x"46", -- 0x08E8
    x"78",x"FE",x"00",x"28",x"0B",x"FE",x"FF",x"C2", -- 0x08F0
    x"54",x"0A",x"79",x"FE",x"F9",x"FA",x"54",x"0A", -- 0x08F8
    x"23",x"4E",x"23",x"46",x"78",x"FE",x"00",x"28", -- 0x0900
    x"0B",x"FE",x"FF",x"C2",x"54",x"0A",x"79",x"FE", -- 0x0908
    x"F9",x"FA",x"54",x"0A",x"2B",x"2B",x"7E",x"FE", -- 0x0910
    x"00",x"CA",x"CA",x"09",x"2B",x"4E",x"23",x"46", -- 0x0918
    x"21",x"08",x"00",x"09",x"7D",x"FD",x"77",x"01", -- 0x0920
    x"DD",x"6E",x"00",x"DD",x"66",x"01",x"11",x"05", -- 0x0928
    x"00",x"19",x"EB",x"1A",x"6F",x"13",x"1A",x"67", -- 0x0930
    x"E5",x"DD",x"6E",x"02",x"DD",x"66",x"03",x"11", -- 0x0938
    x"00",x"00",x"19",x"7E",x"CB",x"27",x"01",x"00", -- 0x0940
    x"00",x"4F",x"E1",x"09",x"7E",x"F6",x"80",x"FD", -- 0x0948
    x"77",x"03",x"C3",x"00",x"0A",x"FD",x"2A",x"06", -- 0x0950
    x"80",x"DD",x"6E",x"02",x"DD",x"66",x"03",x"11", -- 0x0958
    x"01",x"00",x"19",x"4E",x"23",x"46",x"78",x"FE", -- 0x0960
    x"00",x"28",x"0B",x"FE",x"FF",x"C2",x"54",x"0A", -- 0x0968
    x"79",x"FE",x"E1",x"FA",x"54",x"0A",x"23",x"4E", -- 0x0970
    x"23",x"46",x"78",x"FE",x"00",x"28",x"0B",x"FE", -- 0x0978
    x"FF",x"C2",x"54",x"0A",x"79",x"FE",x"E1",x"FA", -- 0x0980
    x"54",x"0A",x"2B",x"2B",x"7E",x"FE",x"00",x"CA", -- 0x0988
    x"CA",x"09",x"2B",x"4E",x"23",x"46",x"21",x"20", -- 0x0990
    x"00",x"09",x"7D",x"FD",x"77",x"01",x"DD",x"6E", -- 0x0998
    x"00",x"DD",x"66",x"01",x"11",x"05",x"00",x"19", -- 0x09A0
    x"EB",x"1A",x"6F",x"13",x"1A",x"67",x"E5",x"DD", -- 0x09A8
    x"6E",x"02",x"DD",x"66",x"03",x"11",x"00",x"00", -- 0x09B0
    x"19",x"7E",x"CB",x"27",x"01",x"00",x"00",x"4F", -- 0x09B8
    x"E1",x"09",x"7E",x"F6",x"80",x"FD",x"77",x"03", -- 0x09C0
    x"18",x"36",x"DD",x"6E",x"02",x"DD",x"66",x"03", -- 0x09C8
    x"11",x"01",x"00",x"19",x"7E",x"FD",x"77",x"01", -- 0x09D0
    x"DD",x"6E",x"00",x"DD",x"66",x"01",x"11",x"05", -- 0x09D8
    x"00",x"19",x"EB",x"1A",x"6F",x"13",x"1A",x"67", -- 0x09E0
    x"E5",x"DD",x"6E",x"02",x"DD",x"66",x"03",x"11", -- 0x09E8
    x"00",x"00",x"19",x"7E",x"CB",x"27",x"01",x"00", -- 0x09F0
    x"00",x"4F",x"E1",x"09",x"7E",x"FD",x"77",x"03", -- 0x09F8
    x"DD",x"6E",x"02",x"DD",x"66",x"03",x"11",x"03", -- 0x0A00
    x"00",x"19",x"7E",x"FD",x"77",x"00",x"DD",x"6E", -- 0x0A08
    x"00",x"DD",x"66",x"01",x"11",x"05",x"00",x"19", -- 0x0A10
    x"EB",x"1A",x"6F",x"13",x"1A",x"67",x"E5",x"DD", -- 0x0A18
    x"6E",x"02",x"DD",x"66",x"03",x"11",x"00",x"00", -- 0x0A20
    x"19",x"7E",x"CB",x"27",x"01",x"00",x"00",x"4F", -- 0x0A28
    x"E1",x"09",x"23",x"7E",x"DD",x"6E",x"00",x"DD", -- 0x0A30
    x"66",x"01",x"11",x"01",x"00",x"19",x"86",x"FD", -- 0x0A38
    x"77",x"02",x"AF",x"16",x"00",x"DD",x"5E",x"04", -- 0x0A40
    x"FD",x"E5",x"E1",x"FD",x"21",x"01",x"00",x"CD", -- 0x0A48
    x"BE",x"1F",x"18",x"32",x"FD",x"E5",x"DD",x"E5", -- 0x0A50
    x"FD",x"E5",x"FD",x"E5",x"AF",x"16",x"00",x"DD", -- 0x0A58
    x"5E",x"04",x"E1",x"FD",x"21",x"01",x"00",x"CD", -- 0x0A60
    x"BB",x"1F",x"3E",x"00",x"FD",x"E1",x"FD",x"77", -- 0x0A68
    x"01",x"3E",x"80",x"FD",x"77",x"03",x"AF",x"16", -- 0x0A70
    x"00",x"DD",x"E1",x"DD",x"5E",x"04",x"E1",x"FD", -- 0x0A78
    x"21",x"01",x"00",x"CD",x"BE",x"1F",x"C9",x"FD", -- 0x0A80
    x"2A",x"06",x"80",x"3A",x"C3",x"73",x"CB",x"4F", -- 0x0A88
    x"20",x"04",x"CB",x"B8",x"18",x"02",x"CB",x"F8", -- 0x0A90
    x"FD",x"70",x"03",x"E5",x"DD",x"66",x"03",x"DD", -- 0x0A98
    x"6E",x"02",x"7E",x"FD",x"77",x"04",x"EE",x"80", -- 0x0AA0
    x"77",x"23",x"5E",x"7B",x"E6",x"07",x"ED",x"44", -- 0x0AA8
    x"C6",x"08",x"FD",x"77",x"01",x"23",x"56",x"CD", -- 0x0AB0
    x"E8",x"07",x"FD",x"73",x"11",x"23",x"5E",x"7B", -- 0x0AB8
    x"E6",x"07",x"FD",x"77",x"00",x"23",x"56",x"CD", -- 0x0AC0
    x"E8",x"07",x"FD",x"73",x"12",x"2A",x"06",x"80", -- 0x0AC8
    x"11",x"13",x"00",x"19",x"FD",x"56",x"12",x"FD", -- 0x0AD0
    x"5E",x"11",x"01",x"03",x"03",x"CD",x"98",x"08", -- 0x0AD8
    x"DD",x"56",x"05",x"DD",x"5E",x"04",x"DD",x"7E", -- 0x0AE0
    x"06",x"DD",x"E1",x"FD",x"2A",x"06",x"80",x"FD", -- 0x0AE8
    x"77",x"05",x"D5",x"2A",x"06",x"80",x"01",x"06", -- 0x0AF0
    x"00",x"09",x"01",x"0B",x"00",x"7A",x"FE",x"70", -- 0x0AF8
    x"30",x"05",x"CD",x"E2",x"1F",x"18",x"03",x"EB", -- 0x0B00
    x"ED",x"B0",x"2A",x"06",x"80",x"11",x"13",x"00", -- 0x0B08
    x"19",x"D9",x"ED",x"5B",x"06",x"80",x"21",x"08", -- 0x0B10
    x"00",x"19",x"EB",x"D9",x"FD",x"2A",x"06",x"80", -- 0x0B18
    x"FD",x"4E",x"05",x"06",x"09",x"7E",x"91",x"FE", -- 0x0B20
    x"12",x"30",x"0E",x"FE",x"09",x"38",x"02",x"D6", -- 0x0B28
    x"09",x"D9",x"6F",x"26",x"00",x"19",x"7E",x"D9", -- 0x0B30
    x"77",x"23",x"10",x"E9",x"D1",x"2A",x"06",x"80", -- 0x0B38
    x"01",x"11",x"00",x"09",x"01",x"0B",x"00",x"7A", -- 0x0B40
    x"FE",x"70",x"30",x"05",x"CD",x"DF",x"1F",x"18", -- 0x0B48
    x"02",x"ED",x"B0",x"DD",x"E5",x"ED",x"5B",x"06", -- 0x0B50
    x"80",x"21",x"13",x"00",x"19",x"EB",x"01",x"14", -- 0x0B58
    x"00",x"09",x"06",x"09",x"1A",x"13",x"D5",x"11", -- 0x0B60
    x"08",x"00",x"19",x"E5",x"5F",x"16",x"00",x"4F", -- 0x0B68
    x"C5",x"3E",x"09",x"90",x"06",x"00",x"D6",x"03", -- 0x0B70
    x"38",x"03",x"04",x"18",x"F9",x"78",x"FD",x"2A", -- 0x0B78
    x"06",x"80",x"FD",x"86",x"12",x"FD",x"CB",x"03", -- 0x0B80
    x"7E",x"FD",x"21",x"01",x"00",x"20",x"29",x"3E", -- 0x0B88
    x"03",x"CD",x"BB",x"1F",x"C1",x"2A",x"06",x"80", -- 0x0B90
    x"C5",x"11",x"84",x"00",x"19",x"59",x"CB",x"3B", -- 0x0B98
    x"CB",x"3B",x"CB",x"3B",x"16",x"00",x"3E",x"09", -- 0x0BA0
    x"90",x"4F",x"06",x"00",x"09",x"FD",x"21",x"01", -- 0x0BA8
    x"00",x"3E",x"04",x"CD",x"BB",x"1F",x"18",x"21", -- 0x0BB0
    x"CB",x"2F",x"CB",x"2F",x"CB",x"2F",x"FE",x"03", -- 0x0BB8
    x"30",x"17",x"57",x"D5",x"E5",x"3E",x"03",x"CD", -- 0x0BC0
    x"BB",x"1F",x"E1",x"11",x"68",x"00",x"19",x"D1", -- 0x0BC8
    x"FD",x"21",x"01",x"00",x"3E",x"04",x"CD",x"BB", -- 0x0BD0
    x"1F",x"C1",x"E1",x"D1",x"10",x"86",x"DD",x"E1", -- 0x0BD8
    x"D9",x"DD",x"56",x"03",x"DD",x"5E",x"02",x"DD", -- 0x0BE0
    x"46",x"05",x"DD",x"4E",x"04",x"D9",x"DD",x"E5", -- 0x0BE8
    x"E1",x"FD",x"2A",x"06",x"80",x"FD",x"7E",x"04", -- 0x0BF0
    x"87",x"4F",x"06",x"00",x"11",x"06",x"00",x"19", -- 0x0BF8
    x"09",x"5E",x"23",x"56",x"2A",x"06",x"80",x"01", -- 0x0C00
    x"7C",x"00",x"09",x"E5",x"C5",x"01",x"05",x"00", -- 0x0C08
    x"7A",x"FE",x"70",x"30",x"05",x"CD",x"E2",x"1F", -- 0x0C10
    x"18",x"03",x"EB",x"ED",x"B0",x"FD",x"2A",x"06", -- 0x0C18
    x"80",x"C1",x"FD",x"09",x"FD",x"7E",x"04",x"FD", -- 0x0C20
    x"2A",x"06",x"80",x"FD",x"77",x"02",x"D1",x"2A", -- 0x0C28
    x"06",x"80",x"01",x"64",x"00",x"09",x"06",x"04", -- 0x0C30
    x"1A",x"DD",x"BE",x"01",x"D5",x"30",x"16",x"D9", -- 0x0C38
    x"87",x"87",x"87",x"6F",x"26",x"00",x"09",x"E5", -- 0x0C40
    x"D9",x"D1",x"EB",x"C5",x"01",x"08",x"00",x"ED", -- 0x0C48
    x"B0",x"C1",x"EB",x"18",x"30",x"DD",x"96",x"01", -- 0x0C50
    x"D9",x"87",x"87",x"87",x"6F",x"26",x"00",x"19", -- 0x0C58
    x"E5",x"D9",x"D1",x"7A",x"FE",x"70",x"30",x"14", -- 0x0C60
    x"C5",x"E5",x"D5",x"01",x"08",x"00",x"CD",x"E2", -- 0x0C68
    x"1F",x"01",x"08",x"00",x"E1",x"09",x"EB",x"E1", -- 0x0C70
    x"09",x"C1",x"18",x"09",x"EB",x"C5",x"01",x"08", -- 0x0C78
    x"00",x"ED",x"B0",x"C1",x"EB",x"D1",x"13",x"10", -- 0x0C80
    x"AF",x"FD",x"2A",x"06",x"80",x"ED",x"5B",x"06", -- 0x0C88
    x"80",x"21",x"1C",x"00",x"19",x"FD",x"4E",x"00", -- 0x0C90
    x"06",x"00",x"09",x"E5",x"DD",x"E1",x"21",x"64", -- 0x0C98
    x"00",x"19",x"E5",x"3E",x"10",x"08",x"E1",x"56", -- 0x0CA0
    x"23",x"E5",x"01",x"0F",x"00",x"09",x"5E",x"EB", -- 0x0CA8
    x"FD",x"46",x"01",x"AF",x"05",x"FA",x"BC",x"0C", -- 0x0CB0
    x"29",x"17",x"18",x"F8",x"5F",x"CD",x"2F",x"0E", -- 0x0CB8
    x"FD",x"7E",x"00",x"3C",x"FD",x"77",x"00",x"FE", -- 0x0CC0
    x"08",x"28",x"04",x"FE",x"10",x"20",x"05",x"01", -- 0x0CC8
    x"10",x"00",x"DD",x"09",x"DD",x"23",x"08",x"3D", -- 0x0CD0
    x"28",x"03",x"08",x"18",x"C9",x"E1",x"FD",x"CB", -- 0x0CD8
    x"03",x"7E",x"20",x"1F",x"2A",x"06",x"80",x"01", -- 0x0CE0
    x"84",x"00",x"09",x"FD",x"56",x"02",x"FD",x"CB", -- 0x0CE8
    x"03",x"4E",x"20",x"04",x"0E",x"0F",x"18",x"02", -- 0x0CF0
    x"0E",x"00",x"06",x"09",x"7E",x"A1",x"B2",x"77", -- 0x0CF8
    x"23",x"10",x"F9",x"FD",x"7E",x"05",x"FD",x"CB", -- 0x0D00
    x"04",x"7E",x"28",x"02",x"C6",x"09",x"4F",x"2A", -- 0x0D08
    x"06",x"80",x"11",x"13",x"00",x"19",x"06",x"09", -- 0x0D10
    x"77",x"3C",x"23",x"10",x"FB",x"FD",x"CB",x"03", -- 0x0D18
    x"7E",x"20",x"73",x"59",x"16",x"00",x"2A",x"06", -- 0x0D20
    x"80",x"01",x"1C",x"00",x"09",x"FD",x"21",x"09", -- 0x0D28
    x"00",x"3E",x"03",x"CD",x"BE",x"1F",x"FD",x"2A", -- 0x0D30
    x"06",x"80",x"2A",x"06",x"80",x"01",x"84",x"00", -- 0x0D38
    x"09",x"DD",x"2A",x"06",x"80",x"01",x"13",x"00", -- 0x0D40
    x"DD",x"09",x"06",x"09",x"DD",x"7E",x"00",x"DD", -- 0x0D48
    x"23",x"CB",x"3F",x"CB",x"3F",x"CB",x"3F",x"5F", -- 0x0D50
    x"16",x"00",x"C5",x"3E",x"09",x"90",x"06",x"00", -- 0x0D58
    x"FE",x"03",x"38",x"05",x"D6",x"03",x"04",x"18", -- 0x0D60
    x"F7",x"FD",x"86",x"11",x"FE",x"20",x"30",x"17", -- 0x0D68
    x"78",x"FD",x"86",x"12",x"FE",x"18",x"30",x"0F", -- 0x0D70
    x"DD",x"E5",x"E5",x"3E",x"04",x"FD",x"21",x"01", -- 0x0D78
    x"00",x"CD",x"BE",x"1F",x"E1",x"DD",x"E1",x"C1", -- 0x0D80
    x"23",x"13",x"05",x"78",x"FE",x"00",x"20",x"BC", -- 0x0D88
    x"FD",x"2A",x"06",x"80",x"18",x"54",x"06",x"00", -- 0x0D90
    x"C5",x"79",x"80",x"80",x"80",x"4F",x"21",x"00", -- 0x0D98
    x"00",x"11",x"18",x"00",x"78",x"3D",x"FA",x"AC", -- 0x0DA0
    x"0D",x"19",x"18",x"F9",x"FD",x"2A",x"06",x"80", -- 0x0DA8
    x"FD",x"7E",x"12",x"80",x"FE",x"18",x"30",x"2B", -- 0x0DB0
    x"CB",x"3F",x"CB",x"3F",x"CB",x"3F",x"57",x"59", -- 0x0DB8
    x"D5",x"01",x"1C",x"00",x"09",x"ED",x"4B",x"06", -- 0x0DC0
    x"80",x"09",x"E5",x"FD",x"21",x"03",x"00",x"3E", -- 0x0DC8
    x"03",x"CD",x"BE",x"1F",x"E1",x"11",x"68",x"00", -- 0x0DD0
    x"19",x"D1",x"FD",x"21",x"03",x"00",x"3E",x"04", -- 0x0DD8
    x"CD",x"BE",x"1F",x"C1",x"04",x"78",x"FE",x"03", -- 0x0DE0
    x"20",x"AE",x"FD",x"2A",x"06",x"80",x"FD",x"46", -- 0x0DE8
    x"06",x"78",x"FE",x"80",x"28",x"21",x"FD",x"4E", -- 0x0DF0
    x"07",x"FD",x"66",x"11",x"FD",x"6E",x"12",x"B7", -- 0x0DF8
    x"ED",x"42",x"28",x"13",x"2A",x"06",x"80",x"11", -- 0x0E00
    x"08",x"00",x"19",x"FD",x"5E",x"06",x"FD",x"56", -- 0x0E08
    x"07",x"01",x"03",x"03",x"CD",x"0B",x"08",x"FD", -- 0x0E10
    x"2A",x"06",x"80",x"2A",x"06",x"80",x"11",x"13", -- 0x0E18
    x"00",x"19",x"FD",x"5E",x"11",x"FD",x"56",x"12", -- 0x0E20
    x"01",x"03",x"03",x"CD",x"0B",x"08",x"C9",x"FD", -- 0x0E28
    x"CB",x"03",x"46",x"20",x"16",x"DD",x"B6",x"00", -- 0x0E30
    x"DD",x"77",x"00",x"7C",x"DD",x"B6",x"08",x"DD", -- 0x0E38
    x"77",x"08",x"7D",x"DD",x"B6",x"10",x"DD",x"77", -- 0x0E40
    x"10",x"18",x"14",x"B7",x"28",x"03",x"DD",x"77", -- 0x0E48
    x"00",x"7C",x"B7",x"28",x"03",x"DD",x"77",x"08", -- 0x0E50
    x"7D",x"B7",x"28",x"03",x"DD",x"77",x"10",x"FD", -- 0x0E58
    x"CB",x"03",x"7E",x"28",x"3C",x"DD",x"E5",x"01", -- 0x0E60
    x"68",x"00",x"DD",x"09",x"FD",x"46",x"02",x"FD", -- 0x0E68
    x"CB",x"03",x"4E",x"20",x"04",x"0E",x"0F",x"18", -- 0x0E70
    x"02",x"0E",x"00",x"7B",x"B7",x"28",x"08",x"DD", -- 0x0E78
    x"7E",x"00",x"A1",x"B0",x"DD",x"77",x"00",x"7C", -- 0x0E80
    x"B7",x"28",x"08",x"DD",x"7E",x"08",x"A1",x"B0", -- 0x0E88
    x"DD",x"77",x"08",x"7D",x"B7",x"28",x"08",x"DD", -- 0x0E90
    x"7E",x"10",x"A1",x"B0",x"DD",x"77",x"10",x"DD", -- 0x0E98
    x"E1",x"C9",x"C5",x"D9",x"DD",x"66",x"03",x"DD", -- 0x0EA0
    x"6E",x"02",x"7E",x"23",x"4E",x"23",x"46",x"23", -- 0x0EA8
    x"5E",x"23",x"56",x"D9",x"87",x"87",x"5F",x"16", -- 0x0EB0
    x"00",x"23",x"19",x"4E",x"23",x"46",x"23",x"5E", -- 0x0EB8
    x"23",x"56",x"60",x"69",x"C1",x"79",x"48",x"CB", -- 0x0EC0
    x"3F",x"CB",x"3F",x"CB",x"3F",x"CB",x"3F",x"47", -- 0x0EC8
    x"C5",x"DD",x"E5",x"E5",x"D5",x"DD",x"6E",x"04", -- 0x0ED0
    x"DD",x"66",x"05",x"DD",x"23",x"DD",x"23",x"23", -- 0x0ED8
    x"23",x"5E",x"23",x"56",x"D5",x"FD",x"E1",x"D1", -- 0x0EE0
    x"E1",x"7E",x"FD",x"CB",x"00",x"7E",x"28",x"02", -- 0x0EE8
    x"CB",x"FF",x"FD",x"77",x"00",x"23",x"1A",x"D9", -- 0x0EF0
    x"6F",x"26",x"00",x"09",x"FD",x"75",x"01",x"FD", -- 0x0EF8
    x"74",x"02",x"D9",x"13",x"1A",x"D9",x"6F",x"26", -- 0x0F00
    x"00",x"19",x"FD",x"75",x"03",x"FD",x"74",x"04", -- 0x0F08
    x"D9",x"13",x"10",x"BF",x"FD",x"E1",x"01",x"04", -- 0x0F10
    x"00",x"FD",x"09",x"D1",x"FD",x"6E",x"00",x"FD", -- 0x0F18
    x"66",x"01",x"FD",x"23",x"FD",x"23",x"E5",x"DD", -- 0x0F20
    x"E1",x"FD",x"E5",x"D5",x"43",x"CD",x"FA",x"1F", -- 0x0F28
    x"D1",x"FD",x"E1",x"15",x"20",x"E6",x"C9",x"2A", -- 0x0F30
    x"D3",x"73",x"CB",x"6E",x"CC",x"49",x"0F",x"CB", -- 0x0F38
    x"66",x"20",x"05",x"23",x"23",x"23",x"18",x"F2", -- 0x0F40
    x"C9",x"E5",x"CB",x"5E",x"28",x"2B",x"CB",x"76", -- 0x0F48
    x"20",x"0D",x"23",x"5E",x"23",x"56",x"1B",x"7B", -- 0x0F50
    x"B2",x"20",x"34",x"E1",x"E5",x"18",x"2C",x"23", -- 0x0F58
    x"5E",x"23",x"56",x"EB",x"5E",x"23",x"56",x"1B", -- 0x0F60
    x"7B",x"B2",x"20",x"23",x"23",x"5E",x"23",x"56", -- 0x0F68
    x"2B",x"2B",x"72",x"2B",x"73",x"E1",x"E5",x"18", -- 0x0F70
    x"12",x"23",x"35",x"20",x"10",x"E1",x"E5",x"CB", -- 0x0F78
    x"76",x"28",x"08",x"23",x"23",x"7E",x"2B",x"77", -- 0x0F80
    x"2B",x"E1",x"E5",x"CB",x"FE",x"E1",x"C9",x"72", -- 0x0F88
    x"2B",x"73",x"18",x"F9",x"02",x"00",x"02",x"00", -- 0x0F90
    x"02",x"00",x"01",x"94",x"0F",x"11",x"BA",x"73", -- 0x0F98
    x"CD",x"98",x"00",x"2A",x"BA",x"73",x"ED",x"5B", -- 0x0FA0
    x"BC",x"73",x"22",x"D3",x"73",x"36",x"30",x"EB", -- 0x0FA8
    x"22",x"D5",x"73",x"C9",x"01",x"00",x"01",x"00", -- 0x0FB0
    x"01",x"B4",x"0F",x"11",x"BE",x"73",x"CD",x"98", -- 0x0FB8
    x"00",x"3A",x"BE",x"73",x"4F",x"2A",x"D3",x"73", -- 0x0FC0
    x"47",x"11",x"03",x"00",x"B7",x"28",x"08",x"CB", -- 0x0FC8
    x"66",x"20",x"6A",x"19",x"0D",x"20",x"F8",x"CB", -- 0x0FD0
    x"6E",x"20",x"62",x"CB",x"EE",x"CB",x"76",x"28", -- 0x0FD8
    x"5C",x"CB",x"5E",x"28",x"58",x"23",x"5E",x"23", -- 0x0FE0
    x"56",x"D5",x"2A",x"D3",x"73",x"E5",x"CB",x"66", -- 0x0FE8
    x"20",x"2E",x"CB",x"6E",x"20",x"23",x"7E",x"E6", -- 0x0FF0
    x"48",x"FE",x"48",x"20",x"1C",x"23",x"23",x"7E", -- 0x0FF8
    x"BA",x"38",x"16",x"20",x"08",x"2B",x"7E",x"BB", -- 0x1000
    x"38",x"0F",x"28",x"31",x"23",x"56",x"2B",x"5E", -- 0x1008
    x"1B",x"1B",x"1B",x"1B",x"73",x"23",x"72",x"18", -- 0x1010
    x"00",x"E1",x"23",x"23",x"23",x"E5",x"18",x"CE", -- 0x1018
    x"06",x"00",x"B7",x"E1",x"D1",x"E5",x"2A",x"D5", -- 0x1020
    x"73",x"ED",x"52",x"4D",x"6B",x"62",x"23",x"23", -- 0x1028
    x"23",x"23",x"ED",x"B0",x"01",x"08",x"00",x"ED", -- 0x1030
    x"42",x"22",x"D5",x"73",x"E1",x"C9",x"02",x"00", -- 0x1038
    x"01",x"00",x"02",x"00",x"01",x"3E",x"10",x"11", -- 0x1040
    x"BF",x"73",x"CD",x"98",x"00",x"2A",x"C0",x"73", -- 0x1048
    x"3A",x"BF",x"73",x"4F",x"EB",x"2A",x"D3",x"73", -- 0x1050
    x"AF",x"47",x"CB",x"6E",x"28",x"3E",x"E5",x"7E", -- 0x1058
    x"E6",x"10",x"F6",x"20",x"77",x"AF",x"B2",x"20", -- 0x1060
    x"0B",x"B1",x"28",x"02",x"CB",x"F6",x"23",x"73", -- 0x1068
    x"23",x"73",x"18",x"42",x"CB",x"DE",x"79",x"B7", -- 0x1070
    x"28",x"1B",x"D5",x"EB",x"2A",x"D5",x"73",x"EB", -- 0x1078
    x"CB",x"F6",x"23",x"73",x"23",x"72",x"EB",x"D1", -- 0x1080
    x"73",x"23",x"72",x"23",x"73",x"23",x"72",x"23", -- 0x1088
    x"22",x"D5",x"73",x"18",x"21",x"23",x"73",x"23", -- 0x1090
    x"72",x"23",x"18",x"1A",x"CB",x"66",x"20",x"06", -- 0x1098
    x"23",x"23",x"23",x"04",x"18",x"B4",x"D5",x"E5", -- 0x10A0
    x"23",x"23",x"23",x"04",x"36",x"30",x"EB",x"E1", -- 0x10A8
    x"CB",x"A6",x"EB",x"D1",x"18",x"A4",x"E1",x"CB", -- 0x10B0
    x"AE",x"78",x"C9",x"01",x"00",x"01",x"00",x"01", -- 0x10B8
    x"BB",x"10",x"11",x"C2",x"73",x"CD",x"98",x"00", -- 0x10C0
    x"3A",x"C2",x"73",x"4F",x"2A",x"D3",x"73",x"47", -- 0x10C8
    x"11",x"03",x"00",x"B7",x"28",x"08",x"CB",x"66", -- 0x10D0
    x"20",x"0C",x"19",x"0D",x"20",x"F8",x"CB",x"6E", -- 0x10D8
    x"20",x"04",x"CB",x"7E",x"20",x"03",x"AF",x"18", -- 0x10E0
    x"0A",x"CB",x"76",x"20",x"02",x"CB",x"EE",x"CB", -- 0x10E8
    x"BE",x"3E",x"01",x"B7",x"C9",x"0F",x"06",x"01", -- 0x10F0
    x"03",x"09",x"00",x"0A",x"0F",x"02",x"0B",x"07", -- 0x10F8
    x"0F",x"05",x"04",x"08",x"0F",x"D3",x"C0",x"AF", -- 0x1100
    x"DD",x"2A",x"08",x"80",x"DD",x"23",x"DD",x"23", -- 0x1108
    x"FD",x"21",x"D7",x"73",x"06",x"0A",x"DD",x"77", -- 0x1110
    x"00",x"DD",x"23",x"FD",x"77",x"00",x"FD",x"23", -- 0x1118
    x"FD",x"77",x"00",x"FD",x"23",x"05",x"20",x"EE", -- 0x1120
    x"32",x"EB",x"73",x"32",x"EC",x"73",x"32",x"EE", -- 0x1128
    x"73",x"32",x"EF",x"73",x"32",x"F0",x"73",x"32", -- 0x1130
    x"F1",x"73",x"C9",x"00",x"C9",x"7C",x"FE",x"00", -- 0x1138
    x"20",x"04",x"DB",x"FC",x"18",x"02",x"DB",x"FF", -- 0x1140
    x"2F",x"C9",x"DB",x"FC",x"2F",x"32",x"EE",x"73", -- 0x1148
    x"DB",x"FF",x"2F",x"32",x"EF",x"73",x"D3",x"80", -- 0x1150
    x"CD",x"3B",x"11",x"DB",x"FC",x"2F",x"32",x"F0", -- 0x1158
    x"73",x"DB",x"FF",x"2F",x"32",x"F1",x"73",x"D3", -- 0x1160
    x"C0",x"C9",x"DB",x"FC",x"21",x"EB",x"73",x"CB", -- 0x1168
    x"67",x"20",x"08",x"CB",x"6F",x"20",x"03",x"35", -- 0x1170
    x"18",x"01",x"34",x"DB",x"FF",x"CB",x"67",x"20", -- 0x1178
    x"09",x"23",x"CB",x"6F",x"20",x"03",x"35",x"18", -- 0x1180
    x"01",x"34",x"C9",x"7D",x"FE",x"01",x"28",x"1A", -- 0x1188
    x"01",x"EB",x"73",x"7C",x"FE",x"00",x"28",x"01", -- 0x1190
    x"03",x"0A",x"5F",x"AF",x"02",x"CD",x"3D",x"11", -- 0x1198
    x"57",x"E6",x"0F",x"6F",x"7A",x"E6",x"40",x"67", -- 0x11A0
    x"18",x"16",x"D3",x"80",x"CD",x"3D",x"11",x"57", -- 0x11A8
    x"D3",x"C0",x"E6",x"0F",x"21",x"F5",x"10",x"06", -- 0x11B0
    x"00",x"4F",x"09",x"6E",x"7A",x"E6",x"40",x"67", -- 0x11B8
    x"C9",x"CD",x"4A",x"11",x"FD",x"21",x"D7",x"73", -- 0x11C0
    x"DD",x"2A",x"08",x"80",x"DD",x"E5",x"DD",x"7E", -- 0x11C8
    x"00",x"CB",x"7F",x"28",x"1E",x"47",x"11",x"02", -- 0x11D0
    x"00",x"DD",x"19",x"E6",x"07",x"28",x"09",x"3A", -- 0x11D8
    x"EE",x"73",x"21",x"EB",x"73",x"CD",x"20",x"12", -- 0x11E0
    x"78",x"E6",x"18",x"28",x"06",x"3A",x"F0",x"73", -- 0x11E8
    x"CD",x"3F",x"12",x"DD",x"E1",x"DD",x"7E",x"01", -- 0x11F0
    x"CB",x"7F",x"28",x"23",x"47",x"11",x"0A",x"00", -- 0x11F8
    x"FD",x"19",x"11",x"07",x"00",x"DD",x"19",x"E6", -- 0x1200
    x"07",x"28",x"09",x"3A",x"EF",x"73",x"21",x"EC", -- 0x1208
    x"73",x"CD",x"20",x"12",x"78",x"E6",x"18",x"28", -- 0x1210
    x"06",x"3A",x"F1",x"73",x"CD",x"3F",x"12",x"C9", -- 0x1218
    x"4F",x"CB",x"48",x"28",x"04",x"CD",x"B9",x"12", -- 0x1220
    x"79",x"CB",x"40",x"28",x"04",x"CD",x"89",x"12", -- 0x1228
    x"79",x"CB",x"50",x"28",x"09",x"7E",x"DD",x"86", -- 0x1230
    x"02",x"DD",x"77",x"02",x"AF",x"77",x"C9",x"4F", -- 0x1238
    x"CB",x"58",x"28",x"04",x"CD",x"E9",x"12",x"79", -- 0x1240
    x"CB",x"60",x"28",x"03",x"CD",x"50",x"12",x"C9", -- 0x1248
    x"C5",x"D5",x"E5",x"E6",x"0F",x"5F",x"FD",x"46", -- 0x1250
    x"08",x"FD",x"7E",x"09",x"FE",x"00",x"20",x"1A", -- 0x1258
    x"7B",x"B8",x"28",x"05",x"FD",x"73",x"08",x"18", -- 0x1260
    x"1C",x"3E",x"01",x"FD",x"77",x"09",x"21",x"F5", -- 0x1268
    x"10",x"16",x"00",x"19",x"7E",x"DD",x"77",x"04", -- 0x1270
    x"18",x"0B",x"7B",x"B8",x"28",x"07",x"FD",x"73", -- 0x1278
    x"08",x"AF",x"FD",x"77",x"09",x"E1",x"D1",x"C1", -- 0x1280
    x"C9",x"C5",x"D5",x"E6",x"40",x"5F",x"FD",x"46", -- 0x1288
    x"00",x"FD",x"7E",x"01",x"FE",x"00",x"20",x"13", -- 0x1290
    x"7B",x"B8",x"28",x"05",x"FD",x"73",x"00",x"18", -- 0x1298
    x"15",x"3E",x"01",x"FD",x"77",x"01",x"DD",x"73", -- 0x12A0
    x"00",x"18",x"0B",x"7B",x"B8",x"28",x"07",x"FD", -- 0x12A8
    x"73",x"00",x"AF",x"FD",x"77",x"01",x"D1",x"C1", -- 0x12B0
    x"C9",x"C5",x"D5",x"E6",x"0F",x"5F",x"FD",x"46", -- 0x12B8
    x"02",x"FD",x"7E",x"03",x"FE",x"00",x"20",x"13", -- 0x12C0
    x"7B",x"B8",x"28",x"05",x"FD",x"73",x"02",x"18", -- 0x12C8
    x"15",x"3E",x"01",x"FD",x"77",x"03",x"DD",x"73", -- 0x12D0
    x"01",x"18",x"0B",x"7B",x"B8",x"28",x"07",x"FD", -- 0x12D8
    x"73",x"02",x"AF",x"FD",x"77",x"03",x"D1",x"C1", -- 0x12E0
    x"C9",x"C5",x"D5",x"E6",x"40",x"5F",x"FD",x"46", -- 0x12E8
    x"06",x"FD",x"7E",x"07",x"FE",x"00",x"20",x"13", -- 0x12F0
    x"7B",x"B8",x"28",x"05",x"FD",x"73",x"06",x"18", -- 0x12F8
    x"15",x"3E",x"01",x"FD",x"77",x"07",x"DD",x"73", -- 0x1300
    x"03",x"18",x"0B",x"7B",x"B8",x"28",x"07",x"FD", -- 0x1308
    x"73",x"06",x"AF",x"FD",x"77",x"07",x"D1",x"C1", -- 0x1310
    x"C9",x"21",x"00",x"00",x"11",x"00",x"40",x"3E", -- 0x1318
    x"00",x"CD",x"D4",x"18",x"CD",x"E9",x"18",x"CD", -- 0x1320
    x"27",x"19",x"21",x"A3",x"18",x"11",x"60",x"00", -- 0x1328
    x"E5",x"D5",x"7E",x"FE",x"FF",x"28",x"1B",x"47", -- 0x1330
    x"04",x"21",x"C3",x"14",x"11",x"08",x"00",x"10", -- 0x1338
    x"15",x"D1",x"D5",x"FD",x"21",x"01",x"00",x"3E", -- 0x1340
    x"03",x"CD",x"BE",x"1F",x"D1",x"E1",x"13",x"23", -- 0x1348
    x"18",x"DE",x"D1",x"E1",x"18",x"03",x"19",x"18", -- 0x1350
    x"E6",x"21",x"4D",x"14",x"11",x"85",x"00",x"FD", -- 0x1358
    x"21",x"16",x"00",x"3E",x"02",x"CD",x"BE",x"1F", -- 0x1360
    x"21",x"63",x"14",x"11",x"A5",x"00",x"FD",x"21", -- 0x1368
    x"16",x"00",x"3E",x"02",x"CD",x"BE",x"1F",x"21", -- 0x1370
    x"C1",x"14",x"11",x"9B",x"00",x"FD",x"21",x"02", -- 0x1378
    x"00",x"3E",x"02",x"CD",x"BE",x"1F",x"21",x"B4", -- 0x1380
    x"14",x"11",x"AA",x"02",x"FD",x"21",x"0D",x"00", -- 0x1388
    x"3E",x"02",x"CD",x"BE",x"1F",x"21",x"3B",x"14", -- 0x1390
    x"11",x"00",x"00",x"3E",x"04",x"FD",x"21",x"12", -- 0x1398
    x"00",x"CD",x"BE",x"1F",x"06",x"01",x"0E",x"C0", -- 0x13A0
    x"CD",x"D9",x"1F",x"21",x"00",x"80",x"7E",x"FE", -- 0x13A8
    x"AA",x"20",x"4C",x"23",x"7E",x"FE",x"55",x"20", -- 0x13B0
    x"46",x"21",x"24",x"80",x"CD",x"46",x"19",x"11", -- 0x13B8
    x"24",x"80",x"21",x"01",x"02",x"CD",x"51",x"19", -- 0x13C0
    x"21",x"24",x"80",x"CD",x"46",x"19",x"23",x"54", -- 0x13C8
    x"5D",x"CD",x"46",x"19",x"21",x"C1",x"01",x"CD", -- 0x13D0
    x"51",x"19",x"21",x"24",x"80",x"CD",x"46",x"19", -- 0x13D8
    x"23",x"CD",x"46",x"19",x"23",x"11",x"AC",x"02", -- 0x13E0
    x"FD",x"21",x"04",x"00",x"3E",x"02",x"CD",x"BE", -- 0x13E8
    x"1F",x"CD",x"68",x"19",x"06",x"01",x"0E",x"80", -- 0x13F0
    x"CD",x"D9",x"1F",x"2A",x"0A",x"80",x"E9",x"21", -- 0x13F8
    x"79",x"14",x"11",x"AA",x"01",x"FD",x"21",x"0D", -- 0x1400
    x"00",x"3E",x"02",x"CD",x"BE",x"1F",x"21",x"86", -- 0x1408
    x"14",x"11",x"E4",x"01",x"FD",x"21",x"1A",x"00", -- 0x1410
    x"3E",x"02",x"CD",x"BE",x"1F",x"21",x"A0",x"14", -- 0x1418
    x"11",x"27",x"02",x"FD",x"21",x"14",x"00",x"3E", -- 0x1420
    x"02",x"CD",x"BE",x"1F",x"21",x"00",x"8A",x"CD", -- 0x1428
    x"6B",x"19",x"06",x"01",x"0E",x"80",x"CD",x"D9", -- 0x1430
    x"1F",x"18",x"FE",x"00",x"00",x"00",x"F0",x"F0", -- 0x1438
    x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"D0", -- 0x1440
    x"80",x"90",x"B0",x"30",x"40",x"60",x"61",x"68", -- 0x1448
    x"69",x"70",x"71",x"78",x"79",x"80",x"81",x"88", -- 0x1450
    x"89",x"64",x"65",x"6C",x"74",x"75",x"7C",x"84", -- 0x1458
    x"85",x"8C",x"8D",x"62",x"63",x"6A",x"6B",x"72", -- 0x1460
    x"73",x"7A",x"7B",x"82",x"83",x"8A",x"8B",x"66", -- 0x1468
    x"67",x"6D",x"76",x"77",x"7D",x"86",x"87",x"8E", -- 0x1470
    x"8F",x"54",x"55",x"52",x"4E",x"20",x"47",x"41", -- 0x1478
    x"4D",x"45",x"20",x"4F",x"46",x"46",x"42",x"45", -- 0x1480
    x"46",x"4F",x"52",x"45",x"20",x"49",x"4E",x"53", -- 0x1488
    x"45",x"52",x"54",x"49",x"4E",x"47",x"20",x"43", -- 0x1490
    x"41",x"52",x"54",x"52",x"49",x"44",x"47",x"45", -- 0x1498
    x"4F",x"52",x"20",x"45",x"58",x"50",x"41",x"4E", -- 0x14A0
    x"53",x"49",x"4F",x"4E",x"20",x"4D",x"4F",x"44", -- 0x14A8
    x"55",x"4C",x"45",x"2E",x"1D",x"20",x"31",x"39", -- 0x14B0
    x"38",x"32",x"20",x"43",x"4F",x"4C",x"45",x"43", -- 0x14B8
    x"4F",x"1E",x"1F",x"00",x"00",x"00",x"00",x"00", -- 0x14C0
    x"00",x"00",x"00",x"3F",x"7F",x"FF",x"FF",x"F3", -- 0x14C8
    x"F3",x"F0",x"F0",x"00",x"80",x"C0",x"C0",x"C0", -- 0x14D0
    x"C0",x"00",x"00",x"3F",x"7F",x"FF",x"FF",x"F3", -- 0x14D8
    x"F3",x"F3",x"F3",x"00",x"80",x"C0",x"C0",x"C0", -- 0x14E0
    x"C0",x"C0",x"C0",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x14E8
    x"F0",x"F0",x"F0",x"FF",x"FF",x"FF",x"F0",x"F0", -- 0x14F0
    x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",x"00",x"00", -- 0x14F8
    x"00",x"00",x"00",x"F1",x"F1",x"F1",x"7B",x"7B", -- 0x1500
    x"7B",x"3F",x"3F",x"E0",x"E0",x"E0",x"C0",x"C0", -- 0x1508
    x"C0",x"80",x"80",x"1F",x"3F",x"7F",x"79",x"78", -- 0x1510
    x"7F",x"7F",x"3F",x"80",x"C0",x"E0",x"E0",x"00", -- 0x1518
    x"80",x"C0",x"E0",x"F3",x"F3",x"FB",x"FB",x"FB", -- 0x1520
    x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",x"C0", -- 0x1528
    x"C0",x"C0",x"C0",x"F3",x"F3",x"FF",x"FF",x"7F", -- 0x1530
    x"3F",x"00",x"00",x"C0",x"C0",x"C0",x"C0",x"80", -- 0x1538
    x"00",x"00",x"00",x"F0",x"F0",x"FF",x"FF",x"FF", -- 0x1540
    x"FF",x"00",x"00",x"00",x"00",x"C0",x"C0",x"C0", -- 0x1548
    x"C0",x"00",x"00",x"3F",x"1F",x"1F",x"1F",x"0E", -- 0x1550
    x"0E",x"00",x"00",x"80",x"00",x"00",x"00",x"00", -- 0x1558
    x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0",x"F0", -- 0x1560
    x"F0",x"00",x"00",x"1F",x"01",x"79",x"7F",x"3F", -- 0x1568
    x"1F",x"00",x"00",x"E0",x"E0",x"E0",x"E0",x"C0", -- 0x1570
    x"80",x"00",x"00",x"FF",x"F7",x"F7",x"F7",x"F3", -- 0x1578
    x"F3",x"00",x"00",x"C0",x"C0",x"C0",x"C0",x"C0", -- 0x1580
    x"C0",x"00",x"00",x"7E",x"81",x"BD",x"A1",x"A1", -- 0x1588
    x"BD",x"81",x"7E",x"1F",x"04",x"04",x"04",x"00", -- 0x1590
    x"00",x"00",x"00",x"44",x"6C",x"54",x"54",x"00", -- 0x1598
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x15A0
    x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20", -- 0x15A8
    x"00",x"20",x"00",x"50",x"50",x"50",x"00",x"00", -- 0x15B0
    x"00",x"00",x"00",x"50",x"50",x"F8",x"50",x"F8", -- 0x15B8
    x"50",x"50",x"00",x"20",x"78",x"A0",x"70",x"28", -- 0x15C0
    x"F0",x"20",x"00",x"C0",x"C8",x"10",x"20",x"40", -- 0x15C8
    x"98",x"18",x"00",x"40",x"A0",x"A0",x"40",x"A8", -- 0x15D0
    x"90",x"68",x"00",x"20",x"20",x"20",x"00",x"00", -- 0x15D8
    x"00",x"00",x"00",x"20",x"40",x"80",x"80",x"80", -- 0x15E0
    x"40",x"20",x"00",x"20",x"10",x"08",x"08",x"08", -- 0x15E8
    x"10",x"20",x"00",x"20",x"A8",x"70",x"20",x"70", -- 0x15F0
    x"A8",x"20",x"00",x"00",x"20",x"20",x"F8",x"20", -- 0x15F8
    x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20", -- 0x1600
    x"20",x"40",x"00",x"00",x"00",x"00",x"F8",x"00", -- 0x1608
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1610
    x"00",x"20",x"00",x"00",x"08",x"10",x"20",x"40", -- 0x1618
    x"80",x"00",x"00",x"70",x"88",x"98",x"A8",x"C8", -- 0x1620
    x"88",x"70",x"00",x"20",x"60",x"20",x"20",x"20", -- 0x1628
    x"20",x"70",x"00",x"70",x"88",x"08",x"30",x"40", -- 0x1630
    x"80",x"F8",x"00",x"F8",x"08",x"10",x"30",x"08", -- 0x1638
    x"88",x"70",x"00",x"10",x"30",x"50",x"90",x"F8", -- 0x1640
    x"10",x"10",x"00",x"F8",x"80",x"F0",x"08",x"08", -- 0x1648
    x"88",x"70",x"00",x"38",x"40",x"80",x"F0",x"88", -- 0x1650
    x"88",x"70",x"00",x"F8",x"08",x"10",x"20",x"40", -- 0x1658
    x"40",x"40",x"00",x"70",x"88",x"88",x"70",x"88", -- 0x1660
    x"88",x"70",x"00",x"70",x"88",x"88",x"78",x"08", -- 0x1668
    x"10",x"E0",x"00",x"00",x"00",x"20",x"00",x"20", -- 0x1670
    x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"20", -- 0x1678
    x"20",x"40",x"00",x"10",x"20",x"40",x"80",x"40", -- 0x1680
    x"20",x"10",x"00",x"00",x"00",x"F8",x"00",x"F8", -- 0x1688
    x"00",x"00",x"00",x"40",x"20",x"10",x"08",x"10", -- 0x1690
    x"20",x"40",x"00",x"70",x"88",x"10",x"20",x"20", -- 0x1698
    x"00",x"20",x"00",x"70",x"88",x"A8",x"B8",x"B0", -- 0x16A0
    x"80",x"78",x"00",x"20",x"50",x"88",x"88",x"F8", -- 0x16A8
    x"88",x"88",x"00",x"F0",x"88",x"88",x"F0",x"88", -- 0x16B0
    x"88",x"F0",x"00",x"70",x"88",x"80",x"80",x"80", -- 0x16B8
    x"88",x"70",x"00",x"F0",x"88",x"88",x"88",x"88", -- 0x16C0
    x"88",x"F0",x"00",x"F8",x"80",x"80",x"F0",x"80", -- 0x16C8
    x"80",x"F8",x"00",x"F8",x"80",x"80",x"F0",x"80", -- 0x16D0
    x"80",x"80",x"00",x"78",x"80",x"80",x"80",x"98", -- 0x16D8
    x"88",x"78",x"00",x"88",x"88",x"88",x"F8",x"88", -- 0x16E0
    x"88",x"88",x"00",x"70",x"20",x"20",x"20",x"20", -- 0x16E8
    x"20",x"70",x"00",x"08",x"08",x"08",x"08",x"08", -- 0x16F0
    x"88",x"70",x"00",x"88",x"90",x"A0",x"C0",x"A0", -- 0x16F8
    x"90",x"88",x"00",x"80",x"80",x"80",x"80",x"80", -- 0x1700
    x"80",x"F8",x"00",x"88",x"D8",x"A8",x"A8",x"88", -- 0x1708
    x"88",x"88",x"00",x"88",x"88",x"C8",x"A8",x"98", -- 0x1710
    x"88",x"88",x"00",x"70",x"88",x"88",x"88",x"88", -- 0x1718
    x"88",x"70",x"00",x"F0",x"88",x"88",x"F0",x"80", -- 0x1720
    x"80",x"80",x"00",x"70",x"88",x"88",x"88",x"A8", -- 0x1728
    x"90",x"68",x"00",x"F0",x"88",x"88",x"F0",x"A0", -- 0x1730
    x"90",x"88",x"00",x"70",x"88",x"80",x"70",x"08", -- 0x1738
    x"88",x"70",x"00",x"F8",x"20",x"20",x"20",x"20", -- 0x1740
    x"20",x"20",x"00",x"88",x"88",x"88",x"88",x"88", -- 0x1748
    x"88",x"70",x"00",x"88",x"88",x"88",x"88",x"88", -- 0x1750
    x"50",x"20",x"00",x"88",x"88",x"88",x"A8",x"A8", -- 0x1758
    x"D8",x"88",x"00",x"88",x"88",x"50",x"20",x"50", -- 0x1760
    x"88",x"88",x"00",x"88",x"88",x"50",x"20",x"20", -- 0x1768
    x"20",x"20",x"00",x"F8",x"08",x"10",x"20",x"40", -- 0x1770
    x"80",x"F8",x"00",x"F8",x"C0",x"C0",x"C0",x"C0", -- 0x1778
    x"C0",x"F8",x"00",x"00",x"80",x"40",x"20",x"10", -- 0x1780
    x"08",x"00",x"00",x"F8",x"18",x"18",x"18",x"18", -- 0x1788
    x"18",x"F8",x"00",x"00",x"00",x"20",x"50",x"88", -- 0x1790
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1798
    x"00",x"00",x"F8",x"40",x"20",x"10",x"00",x"00", -- 0x17A0
    x"00",x"00",x"00",x"00",x"00",x"70",x"88",x"F8", -- 0x17A8
    x"88",x"88",x"00",x"00",x"00",x"F0",x"48",x"70", -- 0x17B0
    x"48",x"F0",x"00",x"00",x"00",x"78",x"80",x"80", -- 0x17B8
    x"80",x"78",x"00",x"00",x"00",x"F0",x"48",x"48", -- 0x17C0
    x"48",x"F0",x"00",x"00",x"00",x"F0",x"80",x"E0", -- 0x17C8
    x"80",x"F0",x"00",x"00",x"00",x"F0",x"80",x"E0", -- 0x17D0
    x"80",x"80",x"00",x"00",x"00",x"78",x"80",x"B8", -- 0x17D8
    x"88",x"70",x"00",x"00",x"00",x"88",x"88",x"F8", -- 0x17E0
    x"88",x"88",x"00",x"00",x"00",x"F8",x"20",x"20", -- 0x17E8
    x"20",x"F8",x"00",x"00",x"00",x"70",x"20",x"20", -- 0x17F0
    x"A0",x"E0",x"00",x"00",x"00",x"90",x"A0",x"C0", -- 0x17F8
    x"A0",x"90",x"00",x"00",x"00",x"80",x"80",x"80", -- 0x1800
    x"80",x"F8",x"00",x"00",x"00",x"88",x"D8",x"A8", -- 0x1808
    x"88",x"88",x"00",x"00",x"00",x"88",x"C8",x"A8", -- 0x1810
    x"98",x"88",x"00",x"00",x"00",x"F8",x"88",x"88", -- 0x1818
    x"88",x"F8",x"00",x"00",x"00",x"F0",x"88",x"F0", -- 0x1820
    x"80",x"80",x"00",x"00",x"00",x"F8",x"88",x"A8", -- 0x1828
    x"90",x"E0",x"00",x"00",x"00",x"F8",x"88",x"F8", -- 0x1830
    x"A0",x"90",x"00",x"00",x"00",x"78",x"80",x"70", -- 0x1838
    x"08",x"F0",x"00",x"00",x"00",x"F8",x"20",x"20", -- 0x1840
    x"20",x"20",x"00",x"00",x"00",x"88",x"88",x"88", -- 0x1848
    x"88",x"70",x"00",x"00",x"00",x"88",x"88",x"90", -- 0x1850
    x"A0",x"40",x"00",x"00",x"00",x"88",x"88",x"A8", -- 0x1858
    x"D8",x"88",x"00",x"00",x"00",x"88",x"60",x"20", -- 0x1860
    x"60",x"88",x"00",x"00",x"00",x"88",x"50",x"20", -- 0x1868
    x"20",x"20",x"00",x"00",x"00",x"F8",x"10",x"20", -- 0x1870
    x"40",x"F8",x"00",x"38",x"40",x"20",x"C0",x"20", -- 0x1878
    x"40",x"38",x"00",x"40",x"20",x"10",x"08",x"10", -- 0x1880
    x"20",x"40",x"00",x"E0",x"10",x"20",x"18",x"20", -- 0x1888
    x"10",x"E0",x"00",x"40",x"A8",x"10",x"00",x"00", -- 0x1890
    x"00",x"00",x"00",x"A8",x"50",x"A8",x"50",x"A8", -- 0x1898
    x"50",x"A8",x"00",x"01",x"02",x"0E",x"0F",x"08", -- 0x18A0
    x"09",x"12",x"13",x"03",x"04",x"0E",x"0F",x"05", -- 0x18A8
    x"14",x"00",x"00",x"05",x"00",x"10",x"11",x"0A", -- 0x18B0
    x"0B",x"15",x"16",x"06",x"07",x"10",x"11",x"05", -- 0x18B8
    x"14",x"00",x"00",x"01",x"02",x"0E",x"0F",x"03", -- 0x18C0
    x"04",x"0E",x"0F",x"03",x"04",x"0E",x"0F",x"0C", -- 0x18C8
    x"0D",x"17",x"18",x"FF",x"4F",x"7D",x"D3",x"BF", -- 0x18D0
    x"7C",x"F6",x"40",x"D3",x"BF",x"79",x"D3",x"BE", -- 0x18D8
    x"1B",x"7A",x"B3",x"20",x"F8",x"CD",x"DC",x"1F", -- 0x18E0
    x"C9",x"06",x"00",x"0E",x"00",x"CD",x"D9",x"1F", -- 0x18E8
    x"06",x"01",x"0E",x"80",x"CD",x"D9",x"1F",x"3E", -- 0x18F0
    x"02",x"21",x"00",x"18",x"CD",x"B8",x"1F",x"3E", -- 0x18F8
    x"04",x"21",x"00",x"20",x"CD",x"B8",x"1F",x"3E", -- 0x1900
    x"03",x"21",x"00",x"00",x"CD",x"B8",x"1F",x"3E", -- 0x1908
    x"00",x"21",x"00",x"1B",x"CD",x"B8",x"1F",x"3E", -- 0x1910
    x"01",x"21",x"00",x"38",x"CD",x"B8",x"1F",x"06", -- 0x1918
    x"07",x"0E",x"00",x"CD",x"D9",x"1F",x"C9",x"21", -- 0x1920
    x"8B",x"15",x"11",x"1D",x"00",x"FD",x"21",x"60", -- 0x1928
    x"00",x"3E",x"03",x"CD",x"BE",x"1F",x"21",x"A3", -- 0x1930
    x"15",x"11",x"00",x"00",x"FD",x"21",x"01",x"00", -- 0x1938
    x"3E",x"03",x"CD",x"BE",x"1F",x"C9",x"01",x"00", -- 0x1940
    x"00",x"7E",x"FE",x"2F",x"C8",x"23",x"03",x"18", -- 0x1948
    x"F8",x"C5",x"FD",x"E1",x"3E",x"20",x"99",x"1F", -- 0x1950
    x"06",x"00",x"4F",x"09",x"44",x"4D",x"62",x"6B", -- 0x1958
    x"50",x"59",x"3E",x"02",x"CD",x"BE",x"1F",x"C9", -- 0x1960
    x"21",x"00",x"17",x"11",x"FF",x"00",x"1B",x"7A", -- 0x1968
    x"B3",x"20",x"FB",x"2B",x"7C",x"B5",x"20",x"F3", -- 0x1970
    x"C9",x"21",x"00",x"00",x"11",x"00",x"40",x"3E", -- 0x1978
    x"00",x"CD",x"82",x"1F",x"CD",x"85",x"1F",x"06", -- 0x1980
    x"0F",x"0E",x"04",x"CD",x"D9",x"1F",x"CD",x"7F", -- 0x1988
    x"1F",x"21",x"7C",x"1A",x"11",x"25",x"00",x"FD", -- 0x1990
    x"21",x"16",x"00",x"3E",x"02",x"CD",x"BE",x"1F", -- 0x1998
    x"21",x"92",x"1A",x"11",x"65",x"00",x"FD",x"21", -- 0x19A0
    x"17",x"00",x"3E",x"02",x"CD",x"BE",x"1F",x"11", -- 0x19A8
    x"C5",x"00",x"CD",x"CA",x"1A",x"11",x"05",x"01", -- 0x19B0
    x"CD",x"CA",x"1A",x"11",x"45",x"01",x"CD",x"CA", -- 0x19B8
    x"1A",x"11",x"85",x"01",x"CD",x"CA",x"1A",x"11", -- 0x19C0
    x"E5",x"01",x"CD",x"CA",x"1A",x"11",x"25",x"02", -- 0x19C8
    x"CD",x"CA",x"1A",x"11",x"65",x"02",x"CD",x"CA", -- 0x19D0
    x"1A",x"11",x"A5",x"02",x"CD",x"CA",x"1A",x"11", -- 0x19D8
    x"05",x"01",x"CD",x"D7",x"1A",x"11",x"45",x"01", -- 0x19E0
    x"CD",x"DC",x"1A",x"11",x"85",x"01",x"CD",x"E1", -- 0x19E8
    x"1A",x"21",x"C2",x"1A",x"11",x"E5",x"01",x"CD", -- 0x19F0
    x"E4",x"1A",x"21",x"C3",x"1A",x"11",x"25",x"02", -- 0x19F8
    x"CD",x"E4",x"1A",x"21",x"C4",x"1A",x"11",x"65", -- 0x1A00
    x"02",x"CD",x"E4",x"1A",x"21",x"C5",x"1A",x"11", -- 0x1A08
    x"A5",x"02",x"CD",x"E4",x"1A",x"11",x"0F",x"01", -- 0x1A10
    x"CD",x"D7",x"1A",x"11",x"4F",x"01",x"CD",x"DC", -- 0x1A18
    x"1A",x"11",x"8F",x"01",x"CD",x"E1",x"1A",x"11", -- 0x1A20
    x"F1",x"01",x"CD",x"EE",x"1A",x"11",x"31",x"02", -- 0x1A28
    x"CD",x"EE",x"1A",x"11",x"71",x"02",x"CD",x"EE", -- 0x1A30
    x"1A",x"11",x"B1",x"02",x"CD",x"EE",x"1A",x"11", -- 0x1A38
    x"2F",x"02",x"CD",x"D7",x"1A",x"11",x"6F",x"02", -- 0x1A40
    x"CD",x"DC",x"1A",x"11",x"AF",x"02",x"CD",x"E1", -- 0x1A48
    x"1A",x"11",x"FB",x"01",x"CD",x"FB",x"1A",x"11", -- 0x1A50
    x"3B",x"02",x"CD",x"FB",x"1A",x"11",x"7B",x"02", -- 0x1A58
    x"CD",x"FB",x"1A",x"11",x"BB",x"02",x"CD",x"FB", -- 0x1A60
    x"1A",x"2A",x"FA",x"73",x"11",x"20",x"00",x"3E", -- 0x1A68
    x"F4",x"CD",x"82",x"1F",x"06",x"01",x"0E",x"C0", -- 0x1A70
    x"CD",x"D9",x"1F",x"C9",x"54",x"4F",x"20",x"53", -- 0x1A78
    x"45",x"4C",x"45",x"43",x"54",x"20",x"47",x"41", -- 0x1A80
    x"4D",x"45",x"20",x"4F",x"50",x"54",x"49",x"4F", -- 0x1A88
    x"4E",x"2C",x"50",x"52",x"45",x"53",x"53",x"20", -- 0x1A90
    x"42",x"55",x"54",x"54",x"4F",x"4E",x"20",x"4F", -- 0x1A98
    x"4E",x"20",x"4B",x"45",x"59",x"50",x"41",x"44", -- 0x1AA0
    x"2E",x"31",x"20",x"3D",x"20",x"53",x"4B",x"49", -- 0x1AA8
    x"4C",x"4C",x"20",x"31",x"2F",x"4F",x"4E",x"45", -- 0x1AB0
    x"20",x"50",x"4C",x"41",x"59",x"45",x"52",x"32", -- 0x1AB8
    x"33",x"34",x"35",x"36",x"37",x"38",x"54",x"57", -- 0x1AC0
    x"4F",x"53",x"21",x"A9",x"1A",x"FD",x"21",x"16", -- 0x1AC8
    x"00",x"3E",x"02",x"CD",x"BE",x"1F",x"C9",x"21", -- 0x1AD0
    x"BF",x"1A",x"18",x"08",x"21",x"C0",x"1A",x"18", -- 0x1AD8
    x"03",x"21",x"C1",x"1A",x"FD",x"21",x"01",x"00", -- 0x1AE0
    x"3E",x"02",x"CD",x"BE",x"1F",x"C9",x"21",x"C6", -- 0x1AE8
    x"1A",x"FD",x"21",x"03",x"00",x"3E",x"02",x"CD", -- 0x1AF0
    x"BE",x"1F",x"C9",x"21",x"C9",x"1A",x"FD",x"21", -- 0x1AF8
    x"01",x"00",x"3E",x"02",x"CD",x"BE",x"1F",x"C9", -- 0x1B00
    x"02",x"00",x"01",x"00",x"02",x"00",x"01",x"08", -- 0x1B08
    x"1B",x"11",x"BA",x"73",x"CD",x"98",x"00",x"3A", -- 0x1B10
    x"BA",x"73",x"2A",x"BB",x"73",x"4F",x"06",x"00", -- 0x1B18
    x"DD",x"21",x"F2",x"73",x"DD",x"09",x"DD",x"09", -- 0x1B20
    x"DD",x"75",x"00",x"DD",x"74",x"01",x"3A",x"C3", -- 0x1B28
    x"73",x"CB",x"4F",x"28",x"27",x"79",x"FE",x"03", -- 0x1B30
    x"28",x"06",x"FE",x"04",x"28",x"10",x"18",x"1C", -- 0x1B38
    x"06",x"04",x"7D",x"B4",x"20",x"04",x"0E",x"03", -- 0x1B40
    x"18",x"28",x"0E",x"07",x"18",x"24",x"06",x"03", -- 0x1B48
    x"7D",x"B4",x"20",x"04",x"0E",x"7F",x"18",x"1A", -- 0x1B50
    x"0E",x"FF",x"18",x"16",x"FD",x"21",x"76",x"1B", -- 0x1B58
    x"FD",x"09",x"FD",x"09",x"FD",x"7E",x"00",x"FD", -- 0x1B60
    x"46",x"01",x"CB",x"3C",x"CB",x"1D",x"3D",x"20", -- 0x1B68
    x"F9",x"4D",x"CD",x"CA",x"1C",x"C9",x"07",x"05", -- 0x1B70
    x"0B",x"06",x"0A",x"02",x"0B",x"04",x"06",x"03", -- 0x1B78
    x"05",x"00",x"01",x"00",x"01",x"00",x"01",x"00", -- 0x1B80
    x"FE",x"FF",x"02",x"00",x"01",x"80",x"1B",x"11", -- 0x1B88
    x"BA",x"73",x"CD",x"98",x"00",x"3A",x"BA",x"73", -- 0x1B90
    x"ED",x"5B",x"BB",x"73",x"FD",x"2A",x"BF",x"73", -- 0x1B98
    x"2A",x"BD",x"73",x"CD",x"AA",x"1B",x"CD",x"3E", -- 0x1BA0
    x"1D",x"C9",x"FD",x"22",x"FE",x"73",x"DD",x"21", -- 0x1BA8
    x"F2",x"73",x"4F",x"06",x"00",x"FE",x"04",x"20", -- 0x1BB0
    x"07",x"3A",x"C3",x"73",x"CB",x"4F",x"28",x"2C", -- 0x1BB8
    x"FD",x"21",x"FF",x"1B",x"FD",x"09",x"FD",x"7E", -- 0x1BC0
    x"00",x"FE",x"00",x"28",x"1F",x"CB",x"23",x"CB", -- 0x1BC8
    x"12",x"3D",x"20",x"F9",x"C5",x"ED",x"4B",x"FE", -- 0x1BD0
    x"73",x"FD",x"7E",x"00",x"FE",x"00",x"28",x"0B", -- 0x1BD8
    x"CB",x"21",x"CB",x"10",x"3D",x"20",x"F9",x"ED", -- 0x1BE0
    x"43",x"FE",x"73",x"C1",x"E5",x"DD",x"09",x"DD", -- 0x1BE8
    x"09",x"DD",x"6E",x"00",x"DD",x"66",x"01",x"19", -- 0x1BF0
    x"EB",x"E1",x"ED",x"4B",x"FE",x"73",x"C9",x"02", -- 0x1BF8
    x"03",x"00",x"03",x"03",x"05",x"00",x"01",x"00", -- 0x1C00
    x"01",x"00",x"01",x"00",x"FE",x"FF",x"02",x"00", -- 0x1C08
    x"01",x"04",x"1C",x"11",x"BA",x"73",x"CD",x"98", -- 0x1C10
    x"00",x"3A",x"BA",x"73",x"ED",x"5B",x"BB",x"73", -- 0x1C18
    x"FD",x"2A",x"BF",x"73",x"2A",x"BD",x"73",x"F5", -- 0x1C20
    x"FE",x"00",x"20",x"22",x"3A",x"C7",x"73",x"FE", -- 0x1C28
    x"01",x"20",x"1B",x"F1",x"E5",x"2A",x"02",x"80", -- 0x1C30
    x"7B",x"CB",x"27",x"CB",x"27",x"5F",x"19",x"EB", -- 0x1C38
    x"FD",x"E5",x"C1",x"79",x"CB",x"27",x"CB",x"27", -- 0x1C40
    x"4F",x"E1",x"ED",x"B0",x"18",x"07",x"F1",x"CD", -- 0x1C48
    x"AA",x"1B",x"CD",x"01",x"1D",x"C9",x"01",x"00", -- 0x1C50
    x"01",x"00",x"01",x"56",x"1C",x"11",x"BA",x"73", -- 0x1C58
    x"CD",x"98",x"00",x"3A",x"BA",x"73",x"47",x"AF", -- 0x1C60
    x"2A",x"04",x"80",x"77",x"23",x"3C",x"B8",x"20", -- 0x1C68
    x"FA",x"C9",x"01",x"00",x"01",x"00",x"01",x"72", -- 0x1C70
    x"1C",x"11",x"BA",x"73",x"CD",x"98",x"00",x"3A", -- 0x1C78
    x"BA",x"73",x"DD",x"2A",x"04",x"80",x"F5",x"FD", -- 0x1C80
    x"21",x"F2",x"73",x"FD",x"5E",x"00",x"FD",x"56", -- 0x1C88
    x"01",x"7B",x"D3",x"BF",x"7A",x"F6",x"40",x"D3", -- 0x1C90
    x"BF",x"F1",x"2A",x"02",x"80",x"DD",x"4E",x"00", -- 0x1C98
    x"DD",x"23",x"06",x"00",x"09",x"09",x"09",x"09", -- 0x1CA0
    x"06",x"04",x"0E",x"BE",x"ED",x"A3",x"00",x"00", -- 0x1CA8
    x"20",x"FA",x"3D",x"20",x"E5",x"C9",x"02",x"00", -- 0x1CB0
    x"01",x"00",x"01",x"00",x"01",x"B6",x"1C",x"11", -- 0x1CB8
    x"BA",x"73",x"CD",x"98",x"00",x"2A",x"BA",x"73", -- 0x1CC0
    x"4C",x"45",x"79",x"D3",x"BF",x"78",x"C6",x"80", -- 0x1CC8
    x"D3",x"BF",x"78",x"FE",x"00",x"20",x"04",x"79", -- 0x1CD0
    x"32",x"C3",x"73",x"78",x"FE",x"01",x"20",x"04", -- 0x1CD8
    x"79",x"32",x"C4",x"73",x"C9",x"03",x"00",x"FE", -- 0x1CE0
    x"FF",x"02",x"00",x"02",x"00",x"01",x"E5",x"1C", -- 0x1CE8
    x"11",x"BA",x"73",x"CD",x"98",x"00",x"2A",x"BA", -- 0x1CF0
    x"73",x"ED",x"5B",x"BC",x"73",x"ED",x"4B",x"BE", -- 0x1CF8
    x"73",x"E5",x"D5",x"E1",x"11",x"00",x"40",x"19", -- 0x1D00
    x"7D",x"D3",x"BF",x"7C",x"D3",x"BF",x"C5",x"D1", -- 0x1D08
    x"E1",x"0E",x"BE",x"43",x"ED",x"A3",x"00",x"00", -- 0x1D10
    x"C2",x"14",x"1D",x"15",x"FA",x"21",x"1D",x"20", -- 0x1D18
    x"F3",x"C9",x"03",x"00",x"FE",x"FF",x"02",x"00", -- 0x1D20
    x"02",x"00",x"01",x"22",x"1D",x"11",x"BA",x"73", -- 0x1D28
    x"CD",x"98",x"00",x"2A",x"BA",x"73",x"ED",x"5B", -- 0x1D30
    x"BC",x"73",x"ED",x"4B",x"BE",x"73",x"7B",x"D3", -- 0x1D38
    x"BF",x"7A",x"D3",x"BF",x"C5",x"D1",x"0E",x"BE", -- 0x1D40
    x"43",x"ED",x"A2",x"00",x"00",x"C2",x"49",x"1D", -- 0x1D48
    x"15",x"FA",x"56",x"1D",x"20",x"F3",x"C9",x"DB", -- 0x1D50
    x"BF",x"C9",x"DD",x"21",x"96",x"1D",x"18",x"10", -- 0x1D58
    x"DD",x"21",x"B7",x"1D",x"18",x"0A",x"DD",x"21", -- 0x1D60
    x"E5",x"1D",x"18",x"04",x"DD",x"21",x"07",x"1E", -- 0x1D68
    x"D9",x"08",x"DD",x"E5",x"08",x"F5",x"08",x"F1", -- 0x1D70
    x"D9",x"D5",x"D9",x"D1",x"FD",x"21",x"01",x"00", -- 0x1D78
    x"2A",x"06",x"80",x"CD",x"A3",x"1B",x"DD",x"E1", -- 0x1D80
    x"DD",x"E5",x"DD",x"E9",x"13",x"0B",x"78",x"B1", -- 0x1D88
    x"D9",x"20",x"E1",x"DD",x"E1",x"C9",x"2A",x"06", -- 0x1D90
    x"80",x"01",x"08",x"00",x"E5",x"D1",x"09",x"EB", -- 0x1D98
    x"CD",x"00",x"1F",x"CD",x"72",x"1E",x"CD",x"5D", -- 0x1DA0
    x"1E",x"FE",x"01",x"20",x"06",x"CD",x"89",x"1E", -- 0x1DA8
    x"CD",x"9A",x"1E",x"D9",x"23",x"18",x"D5",x"2A", -- 0x1DB0
    x"06",x"80",x"01",x"08",x"00",x"E5",x"D1",x"09", -- 0x1DB8
    x"EB",x"CD",x"4E",x"1F",x"CD",x"72",x"1E",x"CD", -- 0x1DC0
    x"5D",x"1E",x"FE",x"01",x"20",x"13",x"CD",x"89", -- 0x1DC8
    x"1E",x"2A",x"06",x"80",x"01",x"08",x"00",x"E5", -- 0x1DD0
    x"D1",x"09",x"EB",x"CD",x"4E",x"1F",x"CD",x"9A", -- 0x1DD8
    x"1E",x"D9",x"23",x"18",x"A7",x"2A",x"06",x"80", -- 0x1DE0
    x"01",x"08",x"00",x"E5",x"D1",x"09",x"EB",x"CD", -- 0x1DE8
    x"12",x"1F",x"CD",x"72",x"1E",x"CD",x"5D",x"1E", -- 0x1DF0
    x"FE",x"01",x"20",x"06",x"CD",x"89",x"1E",x"CD", -- 0x1DF8
    x"9A",x"1E",x"D9",x"23",x"C3",x"8C",x"1D",x"2A", -- 0x1E00
    x"06",x"80",x"01",x"08",x"00",x"E5",x"D1",x"09", -- 0x1E08
    x"EB",x"CD",x"AB",x"1E",x"08",x"F5",x"08",x"F1", -- 0x1E10
    x"D9",x"E5",x"D9",x"D1",x"2A",x"06",x"80",x"01", -- 0x1E18
    x"08",x"00",x"09",x"FD",x"21",x"04",x"00",x"CD", -- 0x1E20
    x"27",x"1C",x"CD",x"5D",x"1E",x"FE",x"01",x"20", -- 0x1E28
    x"24",x"CD",x"89",x"1E",x"2A",x"06",x"80",x"01", -- 0x1E30
    x"08",x"00",x"E5",x"D1",x"09",x"EB",x"CD",x"EA", -- 0x1E38
    x"1E",x"3E",x"04",x"D9",x"E5",x"D9",x"D1",x"2A", -- 0x1E40
    x"06",x"80",x"01",x"08",x"00",x"09",x"FD",x"21", -- 0x1E48
    x"04",x"00",x"CD",x"27",x"1C",x"D9",x"23",x"23", -- 0x1E50
    x"23",x"23",x"C3",x"8C",x"1D",x"08",x"F5",x"08", -- 0x1E58
    x"F1",x"FE",x"03",x"20",x"0A",x"21",x"C3",x"73", -- 0x1E60
    x"CB",x"4E",x"28",x"03",x"3E",x"01",x"C9",x"3E", -- 0x1E68
    x"00",x"C9",x"08",x"F5",x"08",x"F1",x"D9",x"E5", -- 0x1E70
    x"D9",x"D1",x"2A",x"06",x"80",x"01",x"08",x"00", -- 0x1E78
    x"09",x"FD",x"21",x"01",x"00",x"CD",x"27",x"1C", -- 0x1E80
    x"C9",x"3E",x"04",x"D9",x"D5",x"D9",x"D1",x"2A", -- 0x1E88
    x"06",x"80",x"FD",x"21",x"01",x"00",x"CD",x"A3", -- 0x1E90
    x"1B",x"C9",x"3E",x"04",x"D9",x"E5",x"D9",x"D1", -- 0x1E98
    x"2A",x"06",x"80",x"FD",x"21",x"01",x"00",x"CD", -- 0x1EA0
    x"27",x"1C",x"C9",x"E5",x"DD",x"E1",x"D5",x"FD", -- 0x1EA8
    x"E1",x"01",x"08",x"00",x"DD",x"7E",x"00",x"DD", -- 0x1EB0
    x"23",x"57",x"1E",x"04",x"CB",x"17",x"CB",x"14", -- 0x1EB8
    x"CB",x"12",x"CB",x"14",x"1D",x"20",x"F5",x"1E", -- 0x1EC0
    x"04",x"CB",x"17",x"CB",x"15",x"CB",x"12",x"CB", -- 0x1EC8
    x"15",x"1D",x"20",x"F5",x"FD",x"74",x"00",x"FD", -- 0x1ED0
    x"75",x"10",x"FD",x"23",x"FD",x"74",x"00",x"FD", -- 0x1ED8
    x"75",x"10",x"FD",x"23",x"0B",x"79",x"B0",x"20", -- 0x1EE0
    x"CB",x"C9",x"01",x"10",x"00",x"E5",x"7E",x"23", -- 0x1EE8
    x"12",x"13",x"12",x"13",x"0B",x"79",x"FE",x"08", -- 0x1EF0
    x"20",x"01",x"E1",x"79",x"B0",x"20",x"EF",x"C9", -- 0x1EF8
    x"01",x"08",x"00",x"46",x"3E",x"80",x"CB",x"10", -- 0x1F00
    x"1F",x"30",x"FB",x"12",x"23",x"13",x"0D",x"20", -- 0x1F08
    x"F2",x"C9",x"E5",x"DD",x"E1",x"EB",x"01",x"08", -- 0x1F10
    x"00",x"DD",x"CB",x"00",x"16",x"CB",x"1E",x"DD", -- 0x1F18
    x"CB",x"01",x"16",x"CB",x"1E",x"DD",x"CB",x"02", -- 0x1F20
    x"16",x"CB",x"1E",x"DD",x"CB",x"03",x"16",x"CB", -- 0x1F28
    x"1E",x"DD",x"CB",x"04",x"16",x"CB",x"1E",x"DD", -- 0x1F30
    x"CB",x"05",x"16",x"CB",x"1E",x"DD",x"CB",x"06", -- 0x1F38
    x"16",x"CB",x"1E",x"DD",x"CB",x"07",x"16",x"CB", -- 0x1F40
    x"1E",x"23",x"0D",x"20",x"CC",x"C9",x"01",x"07", -- 0x1F48
    x"00",x"09",x"03",x"7E",x"12",x"13",x"2B",x"0B", -- 0x1F50
    x"78",x"B1",x"20",x"F7",x"C9",x"FF",x"FF",x"FF", -- 0x1F58
    x"FF",x"C3",x"00",x"03",x"C3",x"88",x"04",x"C3", -- 0x1F60
    x"C7",x"06",x"C3",x"5A",x"1D",x"C3",x"60",x"1D", -- 0x1F68
    x"C3",x"66",x"1D",x"C3",x"6C",x"1D",x"C3",x"4A", -- 0x1F70
    x"11",x"C3",x"8B",x"11",x"C3",x"79",x"19",x"C3", -- 0x1F78
    x"27",x"19",x"C3",x"D4",x"18",x"C3",x"E9",x"18", -- 0x1F80
    x"C3",x"6A",x"11",x"C3",x"0E",x"1B",x"C3",x"8C", -- 0x1F88
    x"1B",x"C3",x"10",x"1C",x"C3",x"5A",x"1C",x"C3", -- 0x1F90
    x"76",x"1C",x"C3",x"9A",x"0F",x"C3",x"B8",x"0F", -- 0x1F98
    x"C3",x"44",x"10",x"C3",x"BF",x"10",x"C3",x"BC", -- 0x1FA0
    x"1C",x"C3",x"ED",x"1C",x"C3",x"2A",x"1D",x"C3", -- 0x1FA8
    x"55",x"06",x"C3",x"03",x"02",x"C3",x"51",x"02", -- 0x1FB0
    x"C3",x"1D",x"1B",x"C3",x"A3",x"1B",x"C3",x"27", -- 0x1FB8
    x"1C",x"C3",x"66",x"1C",x"C3",x"82",x"1C",x"C3", -- 0x1FC0
    x"AA",x"0F",x"C3",x"C4",x"0F",x"C3",x"53",x"10", -- 0x1FC8
    x"C3",x"CB",x"10",x"C3",x"37",x"0F",x"C3",x"3B", -- 0x1FD0
    x"02",x"C3",x"CA",x"1C",x"C3",x"57",x"1D",x"C3", -- 0x1FD8
    x"01",x"1D",x"C3",x"3E",x"1D",x"C3",x"64",x"06", -- 0x1FE0
    x"C3",x"79",x"06",x"C3",x"C1",x"11",x"C3",x"13", -- 0x1FE8
    x"02",x"C3",x"5E",x"02",x"C3",x"7F",x"02",x"C3", -- 0x1FF0
    x"A3",x"04",x"C3",x"D8",x"06",x"C3",x"3B",x"00"  -- 0x1FF8
  );

begin

	p_rom : process
	begin
		wait until rising_edge(CLK);
		if (ENA = '1') then
			DATA <= ROM(to_integer(unsigned(ADDR)));
		else
			DATA	<= (others => 'Z');
		end if;
	end process;
end RTL;
